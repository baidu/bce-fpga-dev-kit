`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
XcYCcrT1PS/fwGJorpXrEgGilDqsJzT2KK8Nn4QymuGT5XlhqSFqfGeWaEojJw/As0qActVg0S0h
hfpsILZwig==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LqhxCxy/ErdRi+6t8QNU9ARqdr/3bhngsNvmyjYk2DNWNxIiu8yNMUp+HFxCFLGS8UP6dJ0hfyJQ
olpEEz2+fzt3Zae8sW9TrpIghtLZZrTB1WnU+s6Oh1Pib7Kh2sVvKOBgbpVOQ79hLGNYwo/bAjGe
JLIiiXLE6YbygYM2ecg=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GIIb4daF7tXUjQgp+fTa22OSK1LUyaNHxVCcHQ6jwSRe4gjimPQbOcBh8OzQ0fFKWP8qQjj5lJqt
z2cI7aasxAtdQagVpnxCsDyTeZjAk2jqpCW1IZyDxgxX+EI8OgEglrFdUnGJOWZtlH5BEfwGLNXq
OzPvgKGFznoneBMqJHc=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TMBqviXcgKwCBBsPgH8M0zl5GFraJU+H9adhdbX5KtTQs99Um5m5R9I2RZXQw3zgN+ApohHSFJP5
aK2I3/Fmws4LdL9HSYuRJh3t9MH5OV03SNBXRUidIPKA/QWrmxzgOAg+EM5mTNlsdeewmeyn32yq
DadvdXiOD5Sjnhvs2zwIBGh3lDqf4m6M99FdDlad5aAJmsaC5s8MePf/mfhN/yAuBfhZgUGoTGju
LXdCFdOC7MhH5Rr5Lvfm5uq8WaPU7CVPCObbX4uhdDzrHBftl81Wtcq6A07rP82R0rKFTjD8dxKS
kVop+Wm4o3uNxIe6ZZ7FLytVstZQ7PDKT51MKg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YtBxJPKn9np6u3Q1FbxWeViaA0L3GaD1iO44Z+eB+NVSJvlDumqkdY3Zp8bhHAL7PvwuKm8kGEjv
WL+CotdBfypoAahwDr9D5HEyxVBohFrldLPV7dXNwSrB4rEWQyli9mFt34DG+mLyRPDBo4+H06aT
9/ElAoTL2h7MHytPPdc1aItOIVfQEweZkaPGuzaH9Dpc55XL0RQJ5MfnZmdvzF4iwhX2MampY7KJ
Xt6k/QrU8as3c5VEBVDJ4HCZKbvdISqNWFVQzF5Owuq47elXdf4Uid2wVN+PrDJaTP1JVJxAPxEk
kkJViofdygH19HURVLkMqifbY47SUw+CnJf/cQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ma56gNl2N0LNMEI/dU6332/+KOVRvCDFFuJN8oK/IEFguecFg7Xse3lI+Ev9qT6sF8zMNewnvTW1
3TX9iuZxyhBnxoI+En1d0rdpxSzDUZqHXQWoZUMPSRgje053sk4kYfVXiufNQx9DfFocf8ZzRUMA
S2QgGtyncbJ3mU7NsgWZ9M70l+buHoCMmPdmpY+RsOkEJ4L97wx5RCXqEN6B0n1SKSS2Jmnl2XvH
/06FBpWkmT5NDcXNCusfLlJObTN/qZkco9EN5YRMbjZIkL6itQV4V2t7QBY0M43c6mwhhMUg3zFN
uOxqmRbAFDWLbYys0FasRCF7p9TztxbnJ72RRQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
c0G7bSZkmzJzC0ZQnsbJvl4QLvzRPO3aavnGMnfH2+VkFE/XFe7i73LU+3owl1kj+SVeMk00BG3L
6VQbpW2C7bqVjO0aMkntJX6qXjryNEPIqOGeGgYu+WgyVSp9YJ6WkCuMduwOe0FCRXS6hHieq8q3
tiVzLdxFcwva62MRp2oU92nEr62eB3GsCFgrQzsmxoTqlCHI1jAPKI0KLa1A6avkJrpaX611yuDH
zom0MyO8g25fHZSX+pwDEJwZ7OIZAdFvEAsQPMDDu3tTcvVt9tK0uWwGCRovHxBO45Fen5Sv9N8N
jkqy0QzUloIonYB/jpfOh7bZvPjBpDBe+EkiQ9Y4EccTSLnCjjUDPee/cKjjBd2LFCgbVwvg+FOY
tXgdy1u8aIimV3xsTElp6UU3mZTUtFQqbIQwipobSt9TOOevMk23q2wRcejUDvY9X6oEtf2GwX0L
SfOWre0BrkG1gyJZ2O/6BA6LWAfZLgzobns2DA/rf6YlSPyGZtToDvqOaT+YH+ooA0/PFC33fBFb
tsu1fIzMd6PBq3xjzelcddf0xfh+/Hfl/PFD47PZC37150V2rxc4WfdGdd+eNvb0KzyaMBAqamU3
Ppbnrv9j5zhgRBAzUYsLsachuEn8U5NaG8R1YQ89cPu4sd0JmKT4+Xu7trKdOdvkDNZk9bc7VzMM
RHEgyxqwDSqRMjt51X88OacRO5HEMw1qWQmiFvsCYve7PK8HHXx8v+h7wqgc0MQPZh5M0YK6IEyv
59PI7bCctfhX0V8Mn8nor+2ghClIhjfBFG40sB40rSOVniNs9JTAu8hAAawWOqXekcoz6kKsaZUX
SSweLYM0YejlQYttheqnEZxqxKAqZb7c3WYHYCPszNlkmtOj3TsSmwkcmN/MtYiXBvFXawICKOhc
IdQLWWHhlSPjn4YN7jGmKRCozwbu1h64HRVjBZ519Wc1UKxs0DFxAGR5RFjTjHvNHVKJDSuwtLmE
jgM6k77gwXyy/FYqhgdW5aJrveHoED4EGmJFYsaU5jxGgPet1Mm7akXp5UV8KkT5QTTS+RdUuWtU
qGZhc7/LXyBjvBqDewnE6FH4rxC9pJU3q2IxPEnWZWEQGC+VkBlBOgCvOAU1upOUcmrNM3TIj2Pf
m4MdZZr1K/HoumjDoOkLreOKxL5DMjqxnCfD3cua5bKEa+juUVjdt8lQmK+hNYQUJnqkYk9T7zi5
RWlxDiQXs6si4IO6c9qBbuDOwJc4gAfX4RcvvDU55sA2d0uwAvfsrlQCAOGi64HPc5q0oUw5PiOG
YVK46l7sdwpkP5vaUEjrMGFdPm4CivoQMYyV287BTF8dQgi2nXpt14XS25SGWJxA2WVuXE/PF4B6
yVxK8BvLaD5BkdKcKKV3Be04yYfIGREqIIIlIGNb3nVQa56ZLo/KoAZSjuF2f0jWArsPKnwjEWMK
zNUAjGdJEMbhiVJeeO24aSAh+QLFp0Y0f0ESGI/cL/Z3Ycyef3yr9wLAUtZsASmG1/2BtRA5oYrN
CP/hQtAZBw14FM5RSoWwyZmsiYpltvYFXyHkDw2y8HmoCWrVwO/KmW9jzgaoZ1PSCAnIfGtroVMQ
UhZZtRoXLMNFuVfIJO8A1LPfpVfNI+Je+qufy8w7AFwDL7vje4czdJIcN5nYBmFDU3XHc0V1OPSl
14tfiPYDWfIlJV1JX13657PB1KfsQTxh1y66ED2TVml8M5f5hmwOjgcwQW5+/hSTQ4fKOXUS0xDB
xMFicpaKh+r26PewxTFUF2of88uaFOttpba+DxMGMg87rwVnYbqz7Oj94d8tnZ7OVJd7Gb7q32L2
CF4DI1RHU0VlJgdnLKnZIYSboJKOUmyx5/QTr98u8yK0NmmOwfDpxbQW94rqLqpXegV/x9gnOfCs
FtI88wUioUsuy47+2KHX4IbwauJbprXTE10aS3mqNsVXxV53HOmEiwEQQTgg0qixZ96u1PpAUbnt
/J5nDeZzy0knTbDfuPuuNaduqG7WPQgcH7/p5dU+dW2Tlqn2yPCRZA+323JddAYW4UL6OlhsUL+x
A4kOIfctRXNIx2PTFnHBa4ItcYO8aAjRqhCsHzpVy8+w6jBSn8s0YDLx4VT7V7Eq6+TKHVWoop8g
N1fopTciBSi/YNgBQpzbVWriR4PtaZFe5uIBo/LUOvKOOIMRiqfdCK0vzPBUcNwvjOoKgXanaMCt
3vvTPJ4eAIk9YRnBgkB0vBOY0MUn+AP4EupVnAZ625NHXlVSdy+5ciLaYhqpbsFJGuBrNeUnT5Sy
9+kAjH8RndieBA4P2rvdpzNueYwzxJFtaCTELW2mBcgdR32UCfF4dh5AFc2xxC1FE3twant2AgXm
LtRZMO8EUqCIsqQraj8l2BHNlHqId++FTWU62wE/V+jJguNee+b5Y9d5WuA3JoC3Hdu0Fue0AuR/
/fNq8bbBAb7mTdcxil//ep6E1XdZbXNc/s5ckiA2jAYMkX5jUbe6oLfCR3dc6Ysqct/ZKKchtz2G
6QtIX1DZmabhnVVhxmmTaNclIB2A0yxkD38EB04bt/zzFfEqnpFEx31+r+deOdTSjMyFQgydYUfB
pkQyg/1o0/F78b/qqZtpfbzUAdvtq/w8H47t33pZEgtUvs7HXB7ngIXDTQxJR0ycppLl18s3oGm7
BcT55Xo5gGJVbTm7Sa+28AD5mrzwHvH1tjrMmNuGz4h7KpAW01p2q5DvhOi1zBImPMu0JRNBihno
MJIFTfCGkNyVnbW0XmIOKgU+XFrMn7TnbppAN8ygplHOR5ehoP9dTpFt+cuAK6kzTb9zLvAmiu4S
tcuQnwa4/S/93e9UUSYQQ3wenwoVDtm/kUAqEicSo9FJ1IA0jG8bEcTSSfB1rZSbTCXtgrRvSeoF
0kM0wOY/QpEbIeR4GCEctj9+c+PnjNAfHqZX210fz/o2esZJ+43t4IypLfvDM86r+WdzgWpkwqfR
bzJfQifyEFEpfnNgA44Gl0R1fkcQjdJ1S9W1WJmWb0xgjt9fOpP1vv+/KUxjrdtdCOPlbHVR8b4e
opP/j9oUo+u3/iBficjEm3FeE623jQmVhENn/iV0WhmgO/SSpwB+EEuwGGDRWqwrf7eDc89VDWLN
vaci4RxuRiYKZPETZLMslJEJLSxrGUHic8b1/Sk0jtqkTnKaCHokOlApqC2W8X5qnK3oKwpupDbU
2sv4MGNUs2tSrQR2MtALnU/dyptElfljjuScEpBuWvH8SySHeFItSWBiTDJ2egi/B+5Cjw7u7cjX
jEQErkiojpt+MeXh34NVMbocoi7bTYSkM3MiF5Hj8lujo8lpTIkPCpHMuEjul3ww2mlTUIJzDuga
Y75Ra2w43WPfwAFNEKQMMmmLeYC+R3YJH1RkeKodbkT7qmZSsRGDXNGHCmoLLPZA73kE22gPgmtX
pr4M690HCHh6RMqFqJdD7qPJkp62mOUMNigAV1KwGhJ/oG4d43TVB+zcw32rh05TZrxxu3jDdAcG
u3dDhAeq3/ny9Jmeda5oq4ml3K2qBkwOx3m6rg62dQqbMYsK1iyApgUHD2tl4XU6L+3dHVw+4Q0g
Yj+55O0Tl0mXzF3Y+Pm8lRp00XZFGiyJWzX3ChMLdNIcrt4pmlGe8i0KWTiLzNEhRNH5x+gPKosz
8q/P97j6Qh6FK4WXJ8fjcaIzG1BsaGCCcBwRQlyslhSK5Q8+0+aBZSiWqtikinJO3LbGCCVAQlhr
ftfvB3U62y3SPY/KQjMOuTGqFLSBbCekRHGRMEXRSt3LRM8z8DIdA6I2oNAnKdiQlELFGLcaRNTV
chm/LYZRAjY8g/f+9qTNF/12NS/Exy3qK3MzhzQuRQ6mJ5jDY/ETVkgFns9q29CdyrhHB2OkoFF+
o/zylbLf3mfdguoI71Jy85zG7ARd9VcgwSoL4Ortr0a2UGRAU3JNcJeI+OUPwEHZ3xGG29DOxbbg
x5ukuoau4oUG0EGZW+22ioWxiTaX50cJ3E/U3lKZC+AMmpWhCIf8/EzCtSeDu4Vwr5+0cp7ilVyN
hMN7b6YhwQz9D5c/t5z/nGsyipiRBI9Iadmu6XdkkS8/aydNNUkrsn9hnFUSbOxf/aT40h/7y7po
FdUtPrObcS2Zf256twsMGoSAH2aeJvKgxgt/UJKPDoRZ9rDb224cJ8VXkvl0M0CyT7+HMJYEd+z0
dw==
`pragma protect end_protected
