    S_AXI_araddr,
    S_AXI_arburst,
    S_AXI_arcache,
    S_AXI_arid,
    S_AXI_arlen,
    S_AXI_arlock,
    S_AXI_arprot,
    S_AXI_arqos,
    S_AXI_arregion,
    S_AXI_arready,
    S_AXI_arsize,
    S_AXI_arvalid,
    S_AXI_awaddr,
    S_AXI_awburst,
    S_AXI_awcache,
    S_AXI_awid,
    S_AXI_awlen,
    S_AXI_awlock,
    S_AXI_awprot,
    S_AXI_awqos,
    S_AXI_awregion,
    S_AXI_awready,
    S_AXI_awsize,
    S_AXI_awvalid,
    S_AXI_bid,
    S_AXI_bready,
    S_AXI_bresp,
    S_AXI_bvalid,
    S_AXI_rdata,
    S_AXI_rid,
    S_AXI_rlast,
    S_AXI_rready,
    S_AXI_rresp,
    S_AXI_rvalid,
    S_AXI_wdata,
    S_AXI_wlast,
    S_AXI_wready,
    S_AXI_wstrb,
    S_AXI_wvalid,
    S_AXI_LITE_araddr,
    S_AXI_LITE_arprot,
    S_AXI_LITE_arready,
    S_AXI_LITE_arvalid,
    S_AXI_LITE_awaddr,
    S_AXI_LITE_awprot,
    S_AXI_LITE_awready,
    S_AXI_LITE_awvalid,
    S_AXI_LITE_bready,
    S_AXI_LITE_bresp,
    S_AXI_LITE_bvalid,
    S_AXI_LITE_rdata,
    S_AXI_LITE_rready,
    S_AXI_LITE_rresp,
    S_AXI_LITE_rvalid,
    S_AXI_LITE_wdata,
    S_AXI_LITE_wready,
    S_AXI_LITE_wstrb,
    S_AXI_LITE_wvalid,

    C0_DDR4_act_n,
    C0_DDR4_adr,
    C0_DDR4_ba,
    C0_DDR4_bg,
    C0_DDR4_ck_c,
    C0_DDR4_cke,
    C0_DDR4_cs_n,
    C0_DDR4_dm_n,
    C0_DDR4_dq,
    C0_DDR4_dqs_c,
    C0_DDR4_odt,
    C0_DDR4_reset_n,
    C0_SYS_CLK_clk_n,
    C0_SYS_CLK_clk_p,
    C0_DDR4_ck_t,
    C0_DDR4_dqs_t,

    C1_DDR4_act_n,
    C1_DDR4_adr,
    C1_DDR4_ba,
    C1_DDR4_bg,
    C1_DDR4_ck_c,
    C1_DDR4_cke,
    C1_DDR4_cs_n,
    C1_DDR4_dm_n,
    C1_DDR4_dq,
    C1_DDR4_dqs_c,
    C1_DDR4_odt,
    C1_DDR4_reset_n,
    C1_SYS_CLK_clk_n,
    C1_SYS_CLK_clk_p,
    C1_DDR4_ck_t,
    C1_DDR4_dqs_t,

    C2_DDR4_act_n,
    C2_DDR4_adr,
    C2_DDR4_ba,
    C2_DDR4_bg,
    C2_DDR4_ck_c,
    C2_DDR4_cke,
    C2_DDR4_cs_n,
    C2_DDR4_dm_n,
    C2_DDR4_dq,
    C2_DDR4_dqs_c,
    C2_DDR4_odt,
    C2_DDR4_reset_n,
    C2_SYS_CLK_clk_n,
    C2_SYS_CLK_clk_p,
    C2_DDR4_ck_t,
    C2_DDR4_dqs_t,

    C3_DDR4_act_n,
    C3_DDR4_adr,
    C3_DDR4_ba,
    C3_DDR4_bg,
    C3_DDR4_ck_c,
    C3_DDR4_cke,
    C3_DDR4_cs_n,
    C3_DDR4_dm_n,
    C3_DDR4_dq,
    C3_DDR4_dqs_c,
    C3_DDR4_odt,
    C3_DDR4_reset_n,
    C3_SYS_CLK_clk_n,
    C3_SYS_CLK_clk_p,
    C3_DDR4_ck_t,
    C3_DDR4_dqs_t,

    s_axi_aclk,
    pe_clk,
    pe_clk_rst,
    i_soft_rst_n,
    s_axi_aresetn,
    sys_reset,
    usr_irq_ack,
    usr_irq_req,

    // Debug core signals.
    drck,
    shift,
    tdi,
    update,
    sel,
    tdo,
    tms,
    tck,
    runtest,
    reset,
    capture,
    bscanid);

  input [63:0]S_AXI_araddr;
  input [1:0]S_AXI_arburst;
  input [3:0]S_AXI_arcache;
  input [3:0]S_AXI_arid;
  input [7:0]S_AXI_arlen;
  input [0:0]S_AXI_arlock;
  input [2:0]S_AXI_arprot;
  input [3:0]S_AXI_arqos;
  input [3:0]S_AXI_arregion;
  output [0:0]S_AXI_arready;
  input [2:0]S_AXI_arsize;
  input [0:0]S_AXI_arvalid;
  input [63:0]S_AXI_awaddr;
  input [1:0]S_AXI_awburst;
  input [3:0]S_AXI_awcache;
  input [3:0]S_AXI_awid;
  input [7:0]S_AXI_awlen;
  input [0:0]S_AXI_awlock;
  input [2:0]S_AXI_awprot;
  input [3:0]S_AXI_awqos;
  input [3:0]S_AXI_awregion;
  output [0:0]S_AXI_awready;
  input [2:0]S_AXI_awsize;
  input [0:0]S_AXI_awvalid;
  output [3:0]S_AXI_bid;
  input [0:0]S_AXI_bready;
  output [1:0]S_AXI_bresp;
  output [0:0]S_AXI_bvalid;
  output [255:0]S_AXI_rdata;
  output [3:0]S_AXI_rid;
  output [0:0]S_AXI_rlast;
  input [0:0]S_AXI_rready;
  output [1:0]S_AXI_rresp;
  output [0:0]S_AXI_rvalid;
  input [255:0]S_AXI_wdata;
  input [0:0]S_AXI_wlast;
  output [0:0]S_AXI_wready;
  input [31:0]S_AXI_wstrb;
  input [0:0]S_AXI_wvalid;
  input [15:0]S_AXI_LITE_araddr;
  input [2:0]S_AXI_LITE_arprot;
  output S_AXI_LITE_arready;
  input S_AXI_LITE_arvalid;
  input [15:0]S_AXI_LITE_awaddr;
  input [2:0]S_AXI_LITE_awprot;
  output S_AXI_LITE_awready;
  input S_AXI_LITE_awvalid;
  input S_AXI_LITE_bready;
  output [1:0]S_AXI_LITE_bresp;
  output S_AXI_LITE_bvalid;
  output [31:0]S_AXI_LITE_rdata;
  input S_AXI_LITE_rready;
  output [1:0]S_AXI_LITE_rresp;
  output S_AXI_LITE_rvalid;
  input [31:0]S_AXI_LITE_wdata;
  output S_AXI_LITE_wready;
  input [3:0]S_AXI_LITE_wstrb;
  input S_AXI_LITE_wvalid;

  output C0_DDR4_act_n;
  output [16:0]C0_DDR4_adr;
  output [1:0]C0_DDR4_ba;
  output [0:0]C0_DDR4_bg;
  output [0:0]C0_DDR4_ck_c;
  output [0:0]C0_DDR4_cke;
  output [0:0]C0_DDR4_cs_n;
  inout [8:0]C0_DDR4_dm_n;
  inout [71:0]C0_DDR4_dq;
  inout [8:0]C0_DDR4_dqs_c;
  output [0:0]C0_DDR4_odt;
  output C0_DDR4_reset_n;
  input C0_SYS_CLK_clk_n;
  input C0_SYS_CLK_clk_p;
  output [0:0]C0_DDR4_ck_t;
  inout [8:0]C0_DDR4_dqs_t;

  output C1_DDR4_act_n;
  output [16:0]C1_DDR4_adr;
  output [1:0]C1_DDR4_ba;
  output [0:0]C1_DDR4_bg;
  output [0:0]C1_DDR4_ck_c;
  output [0:0]C1_DDR4_cke;
  output [0:0]C1_DDR4_cs_n;
  inout [8:0]C1_DDR4_dm_n;
  inout [71:0]C1_DDR4_dq;
  inout [8:0]C1_DDR4_dqs_c;
  output [0:0]C1_DDR4_odt;
  output C1_DDR4_reset_n;
  input C1_SYS_CLK_clk_n;
  input C1_SYS_CLK_clk_p;
  output [0:0]C1_DDR4_ck_t;
  inout [8:0]C1_DDR4_dqs_t;

  output C2_DDR4_act_n;
  output [16:0]C2_DDR4_adr;
  output [1:0]C2_DDR4_ba;
  output [0:0]C2_DDR4_bg;
  output [0:0]C2_DDR4_ck_c;
  output [0:0]C2_DDR4_cke;
  output [0:0]C2_DDR4_cs_n;
  inout [8:0]C2_DDR4_dm_n;
  inout [71:0]C2_DDR4_dq;
  inout [8:0]C2_DDR4_dqs_c;
  output [0:0]C2_DDR4_odt;
  output C2_DDR4_reset_n;
  input C2_SYS_CLK_clk_n;
  input C2_SYS_CLK_clk_p;
  output [0:0]C2_DDR4_ck_t;
  inout [8:0]C2_DDR4_dqs_t;

  output C3_DDR4_act_n;
  output [16:0]C3_DDR4_adr;
  output [1:0]C3_DDR4_ba;
  output [0:0]C3_DDR4_bg;
  output [0:0]C3_DDR4_ck_c;
  output [0:0]C3_DDR4_cke;
  output [0:0]C3_DDR4_cs_n;
  inout [8:0]C3_DDR4_dm_n;
  inout [71:0]C3_DDR4_dq;
  inout [8:0]C3_DDR4_dqs_c;
  output [0:0]C3_DDR4_odt;
  output C3_DDR4_reset_n;
  input C3_SYS_CLK_clk_n;
  input C3_SYS_CLK_clk_p;
  output [0:0]C3_DDR4_ck_t;
  inout [8:0]C3_DDR4_dqs_t;

  input s_axi_aclk;
  input s_axi_aresetn;
  
  input pe_clk;
  input pe_clk_rst;
  input i_soft_rst_n;
  input sys_reset;
  input [15:0]usr_irq_ack;
  output [15:0]usr_irq_req;

  // Debug core signals.
  input  drck;
  input  shift;
  input  tdi;
  input  update;
  input  sel;
  output  tdo;
  input  tms;
  input  tck;
  input  runtest;
  input  reset;
  input  capture;
  output  [31 : 0] bscanid;

  wire [63:0]S_AXI_araddr;
  wire [1:0]S_AXI_arburst;
  wire [3:0]S_AXI_arcache;
  wire [3:0]S_AXI_arid;
  wire [7:0]S_AXI_arlen;
  wire [0:0]S_AXI_arlock;
  wire [2:0]S_AXI_arprot;
  wire [3:0]S_AXI_arqos;
  wire [3:0]S_AXI_arregion;
  wire [0:0]S_AXI_arready;
  wire [2:0]S_AXI_arsize;
  wire [0:0]S_AXI_arvalid;
  wire [63:0]S_AXI_awaddr;
  wire [1:0]S_AXI_awburst;
  wire [3:0]S_AXI_awcache;
  wire [3:0]S_AXI_awid;
  wire [7:0]S_AXI_awlen;
  wire [0:0]S_AXI_awlock;
  wire [2:0]S_AXI_awprot;
  wire [3:0]S_AXI_awqos;
  wire [3:0]S_AXI_awregion;
  wire [0:0]S_AXI_awready;
  wire [2:0]S_AXI_awsize;
  wire [0:0]S_AXI_awvalid;
  wire [3:0]S_AXI_bid;
  wire [0:0]S_AXI_bready;
  wire [1:0]S_AXI_bresp;
  wire [0:0]S_AXI_bvalid;
  wire [255:0]S_AXI_rdata;
  wire [3:0]S_AXI_rid;
  wire [0:0]S_AXI_rlast;
  wire [0:0]S_AXI_rready;
  wire [1:0]S_AXI_rresp;
  wire [0:0]S_AXI_rvalid;
  wire [255:0]S_AXI_wdata;
  wire [0:0]S_AXI_wlast;
  wire [0:0]S_AXI_wready;
  wire [31:0]S_AXI_wstrb;
  wire [0:0]S_AXI_wvalid;
  wire [15:0]S_AXI_LITE_araddr;
  wire [2:0]S_AXI_LITE_arprot;
  wire S_AXI_LITE_arready;
  wire S_AXI_LITE_arvalid;
  wire [15:0]S_AXI_LITE_awaddr;
  wire [2:0]S_AXI_LITE_awprot;
  wire S_AXI_LITE_awready;
  wire S_AXI_LITE_awvalid;
  wire S_AXI_LITE_bready;
  wire [1:0]S_AXI_LITE_bresp;
  wire S_AXI_LITE_bvalid;
  wire [31:0]S_AXI_LITE_rdata;
  wire S_AXI_LITE_rready;
  wire [1:0]S_AXI_LITE_rresp;
  wire S_AXI_LITE_rvalid;
  wire [31:0]S_AXI_LITE_wdata;
  wire S_AXI_LITE_wready;
  wire [3:0]S_AXI_LITE_wstrb;
  wire S_AXI_LITE_wvalid;

  wire s_axi_aclk;
  wire s_axi_aresetn;
  wire pe_clk;
  wire pe_clk_rst;
  wire i_soft_rst_n;
  wire sys_reset;
  wire [15:0]usr_irq_ack;
  wire [15:0]usr_irq_req;

  wire C0_DDR4_act_n;
  wire [16:0]C0_DDR4_adr;
  wire [1:0]C0_DDR4_ba;
  wire [0:0]C0_DDR4_bg;
  wire [0:0]C0_DDR4_ck_c;
  wire [0:0]C0_DDR4_cke;
  wire [0:0]C0_DDR4_cs_n;
  wire [8:0]C0_DDR4_dm_n;
  wire [71:0]C0_DDR4_dq;
  wire [8:0]C0_DDR4_dqs_c;
  wire [0:0]C0_DDR4_odt;
  wire C0_DDR4_reset_n;
  wire C0_SYS_CLK_clk_n;
  wire C0_SYS_CLK_clk_p;
  wire [0:0]C0_DDR4_ck_t;
  wire [8:0]C0_DDR4_dqs_t;

  wire C1_DDR4_act_n;
  wire [16:0]C1_DDR4_adr;
  wire [1:0]C1_DDR4_ba;
  wire [0:0]C1_DDR4_bg;
  wire [0:0]C1_DDR4_ck_c;
  wire [0:0]C1_DDR4_cke;
  wire [0:0]C1_DDR4_cs_n;
  wire [8:0]C1_DDR4_dm_n;
  wire [71:0]C1_DDR4_dq;
  wire [8:0]C1_DDR4_dqs_c;
  wire [0:0]C1_DDR4_odt;
  wire C1_DDR4_reset_n;
  wire C1_SYS_CLK_clk_n;
  wire C1_SYS_CLK_clk_p;
  wire [0:0]C1_DDR4_ck_t;
  wire [8:0]C1_DDR4_dqs_t;

  wire C2_DDR4_act_n;
  wire [16:0]C2_DDR4_adr;
  wire [1:0]C2_DDR4_ba;
  wire [0:0]C2_DDR4_bg;
  wire [0:0]C2_DDR4_ck_c;
  wire [0:0]C2_DDR4_cke;
  wire [0:0]C2_DDR4_cs_n;
  wire [8:0]C2_DDR4_dm_n;
  wire [71:0]C2_DDR4_dq;
  wire [8:0]C2_DDR4_dqs_c;
  wire [0:0]C2_DDR4_odt;
  wire C2_DDR4_reset_n;
  wire C2_SYS_CLK_clk_n;
  wire C2_SYS_CLK_clk_p;
  wire [0:0]C2_DDR4_ck_t;
  wire [8:0]C2_DDR4_dqs_t;

  wire C3_DDR4_act_n;
  wire [16:0]C3_DDR4_adr;
  wire [1:0]C3_DDR4_ba;
  wire [0:0]C3_DDR4_bg;
  wire [0:0]C3_DDR4_ck_c;
  wire [0:0]C3_DDR4_cke;
  wire [0:0]C3_DDR4_cs_n;
  wire [8:0]C3_DDR4_dm_n;
  wire [71:0]C3_DDR4_dq;
  wire [8:0]C3_DDR4_dqs_c;
  wire [0:0]C3_DDR4_odt;
  wire C3_DDR4_reset_n;
  wire C3_SYS_CLK_clk_n;
  wire C3_SYS_CLK_clk_p;
  wire [0:0]C3_DDR4_ck_t;
  wire [8:0]C3_DDR4_dqs_t;

  // Debug core signals.
  wire drck;
  wire shift;
  wire tdi;
  wire update;
  wire sel;
  wire tdo;
  wire tms;
  wire tck;
  wire runtest;
  wire reset;
  wire capture;
  wire [31 : 0] bscanid;
