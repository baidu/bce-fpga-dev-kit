`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
BHK9i0N/ZGXXNgTHeO5ITBPMNfTXpW9yQfuE2YIP4CL8fawovNmbXnJ09yr4zDTR7aw8or1/OSu8
iu8fyVyERA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
THuQBz9qqp70ESgcgwkoYoCncKelGtAG7+/Mp0cX7zI/cxLTh4Pc3yg4X4DZ/Lr0GKKRFtfZ172T
wJ5a+w8AGp9ELO1rVdiPANLr4r2ujaMUlyrCQkwdsZJw9vGHDu3EBmnedTkQ/xUrCLa8yh18fF0U
qt4jPG10LVAnkAkhHtY=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FcHoX+ft6pdL/MbDYWZQYR5rs3rM8KovkmVa/1uQfEA8rlE14ROodRrSkG0BLHroINHLSNsI0M2Z
qrHu3IRiPNkLoKaXEVg1m18nkHRe07f7DMPcBVug9GtaSyh+YfDXM6R7NJV/tw+/aBGzMPl3YPZA
5bZfiErboVNh4sYJI8s=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TliMKvv5uxhWrClZCCZzIc6mhkF9oy15XaC3rX4Eg3juny/DEd1AQgIYv2K4BMqu5aGI8EGyMeeX
ePv5NGX90b3YvXnduyekCw/sEBpl8wbwP1jkAuCoQaFUrIIaOPeDAbr+Z4V0Bit/XGoPmyPYh5Iv
MBzxPiBvt/DdCb5Liw/U70Xkrdz7oQUNsIuZKmPNfhKWjgMyrUu9X+sFRxvmctCTyIu9RzLlLa7/
mKbwVQXEPm8z9n5I83mV5k/hJHNlRlvAVwL0gSlMk1FL84EKemQWJWAUquT9CuR06GSqOF9chAEv
K5WXLva/d/v95pqP7OHFGisYMsrVpQPaJ4SNIA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
D3IYhEzSAAZQuOdBKHRi+1Y4LiiSGJ2TAkNt11HzbjiBzHrGOY7UaUGOUrS39xyqA9wm7TQMqM1J
GyECVN9Vgwzb1JguPDqKM0SQaaTsIUiQ2mx9yK0ugWfTGukh0uznC9TlHHZ/PQ+g33QYR1ZNou2p
IBnsb2ICjpGIGIeBK4zB/ZbJpvL//b20Bd4oPly4UZT0H9SbetVfvTeQHxfpysVbrOQh0z3bWJl0
XvO4OVapKQnfdb9GnAnzrPU+DUjt8T4svBs1pD4ZS+fPGndmzoc4eDxop8dakd/8ymCxCRHRxHvw
7to/KwY2tuPoPBEbA4CR6sS+7oE47wAHF7dRgA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
N4he4pACOUEjAoQxqAX8P6ETlIdtA0OpfiKcoW6XwNSmucCQ8V94DRq075gc6sykeJ3wcFykL1Yo
OAB/fiQ+8B/a34Z15OgiWI35le0kNIpbsc9SvRonXzyDF3WZuUeKWvcNA8t1NkSBcwLPPO9b8zCv
ydobmixV++ivs1BdAiT+8Xmi+Zs7mWzmI7bCX9Sg3/lJe/nnsblyZF6boyk9QFeKCNUUnIxK+vk2
Iz9yQVhkj/88U2PMX/21dzSBnmQCkP8TWLPdlrdpC7GJZ7NK3nFFpXJ85A8+PmDp1EKIx4Wnrc8B
NPoTyrQ8VJPhUv5P5FJsHIz9Ke4RY1UJXmadYw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135936)
`pragma protect data_block
LD+C+SZJfba21h/hbxKPfXDHXyDqUc3joTI85PMnoguUo10Lgn7oYWg2oNQxaLDJbXkZP7vyu17F
jwrLv207zXTXSJB7mR2G5Oz+fpXc8zq5IE3ZQNE5bSRSPh2rgnE/ZSR2+Z2m53PtI1jIAbtcjKks
qdHmcxX30K7j6ZxbncMGhxUiTePIq2QEXpdNNB7j69PaaTQxF0tdMSfMI9pCVsf4hj+c4OHlFwJc
v65yrpHLsqPR7aejm6Bu3I6g6UPmzTQQi4IuIWEbySCgKQ6nqY3Q9yLqxPHjNxzIEFnGD1dQtj6u
2dBZXcwESrkWznhKW7KolFj4J0RaNhLRcNtxmaIsAejy5kwuDJH230xXLJgZ1/ajq0LZ7kXI5MCm
MMtcrdmNlDAlqgZIFT+jMivEMnfAtf3+oMHyDOwxIWGAh09gQEak7q7gjDcxMeMRQlLk7azfjbAC
QHkgGctsdZdyNl3Hx6SOsrlp/BEZn/ghJk6JEJ7tq/22GHyuEFa0EIh51fHhXDQAlSAae3OhLToy
gj8eYCwcFKmCRV0N/e7BexgRAGXG+gM3NkjnDkpBeoo1woeQpxgkDfICzdalZ2XWgKPbhw3qU79G
jaGSCarWnFJ+nUAqLIcP7pRZxQ9Rn9VP25dAn+FG8EmPl14xWMr2dABpHkixSlF40O5aw6v6qcLm
Hbk65la6DqvZqCKR32Gxpmz7Gg1lfooSrC31SweSLMjp4E4e89equImK+JZW/IS45AzlOouNUq4x
0mCKokiR+iouEDP+yltdP2S7sHWFIWj5NrPD+stKaFxD5XCisGdzZdyYEvcwNhs7Ooyajke3Jxty
AL8ddT9a4Xxp9C2Ud5RAaj/t+wxtLV7ckQ+ppqUMiGcaI2roV1JCr15grN7kQZEI+H3jDXOzIuEP
FG3+ZYyWt41yelfZ2lGsGSVRGPy/YIqH+ZrAZNB7+p7zlHceKsfJuAu8KApRYgv5qYTLIvhGbd4s
CuRFUrKwWPEmXP+3koPfK3OaLqya8AA6homzw1rRQ7tTOU733aLesDzv1Brz8DH+w0+S9f9s1gFC
MUi8lPMjqK1l+OHpiO5XpsFTBE8aA/8VVpuG+ZAxfJsVYfsCtv4CNxmEhisSWq2FyLWNoqVnPDhB
eUHGluGwDyiXYk7nxZ4Qsd3XOJAjV0lK6YY0B8EVzTl4kXS4/esOHZHaH//XxHk+/8IxYrbVBqSe
tcPxCcdr87zlFlQV1D/w+XOFO1EFDAz5UZQRGi5rs8Mqx1qx479S5yOJ1fjTwHAc5yRVgGz4e73I
WyLnQH2GO8vGHV3Woya6ghX50Bi2EtYqOhkYSUIb6fUKXpfHbP8bT54KoXmxZq4VbMFGACjU1Lkk
TO9gvAhov/7Dh7mVY2/oFqUE1GAaicX08Nwt0NtkfCAFISRn2g33ecKzNz+ucN5RRDliVRSPAZXH
pFhjdrlSdDelpz4ll9r5HPrU34h8Ono31qQWVcX+oHNKt9IJ5BfbCHWQVzRGPtT9B6NMpq+rYVEE
tP2UJXUYDENtOIv0C23pyrOe5jF87CJu2MIWm1To3TDOw0iyCFOT/vTXWNzOYWmtQnbJnmLG5f4G
n2jAAUxjiRD5BLeOM8w2Trc9ECRGYU7XyZC9R59eXVDGyIJNYehURXqvTRRm5DmSTwQ5CzgkYuoW
ZIjLPYtTF+TnCQAeEp0W2tCpyt34AJaVS5poAW+uE76qci2bBE3OTbU0f3XW78oJ6ekwSw9cKu45
wvsR2LFl92TN1uHU9epzoP64UiQxhN8oM3anCOjBsQcHdgcKRVmXr0tMRKS1vd9rrB8gNHzxc38m
6oFzIDrVgI4CC+1R8TpjWvPfysC6hctGg3hyuPl88bCmb/88UeAEKIIz/fgdpuDxQKE7TinDQMzF
lXgM8YuVXAFYfPlsVPNdzr4b8aO5bJUPjJfkXiqgQeUvqRnErt2EW/x/sQvl9UUThOU+9R5ffmjr
Ma9Ot0km0j49WWs4ogzVCPGvCWCpIfvrdipwEXfoT8AnfQAfYOnexOQh95qq2jTUjDYDplJ4Gc6B
ouB5YkSDCnm19AQIm5VT8rrlfK6ZP1raj0TJD+acExenIRBlxEPe9kdmKiFRHcZYmTjwOa37HLwN
nBO30GJAoerwxpgJ8KxIctzn/CptPwILiM1iQo6aBjrq0TpRgtij47ouUbn5XdGiWa3DwbW0swVm
J3gjlxp4t6ETSdJUCkeZOHn7cTPQ1A90E4cRlo0w4ZhxOUQxbWzaQ1It8NpKV/MtuMT9IijqgAMU
Z8tMCLqO5S9REaGqEFGEcz9WEPRE1Uy02c1JNn9DcvKWRVI9qlFO9YqoxjPOk+2ddAW9ueGb9Wbe
+KNXAO7o4aXCUH4SPsf7x6FSywniqmA5vsP61Q+BQ9oICZR4qgkAKlhAcDnKmc9uvozh4+Lq/1VR
igJgdwuIIGPhr13AX+zCwe2SItEAf3VouMy/0kh2vWjtnCXpeMWW42CKpr772JrR1V5tqNsBMYUA
jlQVpNaWgWBkTv7KCp3WxBtm2Xd9b7rVsC5ZhTGEeh7c3UBflF31FggHcfQVXTYwai6fI2p1A55/
APwmtNO1V2z9XsVssx0PD6/62OYJhg+eXRSHHS3UzbWkVbvhwCv9iyEqhaALxVZ+7hB1DfmM8EaD
ZDsxFxg784Wn7USegTMk8qrygVIe1VhxZbmJmsU9ujiHLBijfWlD1VYlQdUVc1Uq7aQVyJwx/02k
qOgDtjnLLq0AqqfHE9NiU/Qsf0EzYLM1rl78453ccX1ip981SAvIxayHjMtt9DYmJ5lvrQ5dtHOk
X2X2YgGFXxH6Jc7LyjFw3r062LgQy+1iSJi7RS/jKu0NwqGPkxUWbxU9Qmq3ZWRgnO1eeD53GKkh
uBMB8PmHwsNwjcAeM8Z0T9PRsIghxAmMFmXYI2Zvh+l/5DhYPcoX6Jjt+Ibwv9VIt5ym7QXM9+Ee
66Pj79II4yzmeGxClad5lFRHujnN0NkxIpryU4T9kVkvkur/8PdsnyAU9/6EBt4RSCt1TZV99ZP2
JyL0B5PgUF0bm2g2dESjZ9Sde8uBXCu1PeQNRlspmY00rW02OzHCF0vMN6TfQYgjANx1tUXgUWhk
Ius6yfUS2Em79gH2c85UIx9VX01prhsEqfdIjQi9NqOyKkRwbDJUKmId2QlM2Y6aN9LzGsVo3MoX
T1VwaTstvanBmGxWA4/ZpuuHgKY/95nIIg0FA98XDy944Iqgv826BnccicsxjjhzSiwERaGM3rlO
xtW8Gijplqj35hstSzD/jwcW6sqk43whT+1Q+48qndtDTAefByiVgJxH5aZ4/JU6HRhiXKdDns6m
xigtFepUbWA/Ema46cwWT9ncRtHK4Kg/821NtQTntRrGdpzSjDmeedcLINxy1v4ERUosMWw+LBTA
sXUriKje10s6AspJWz5wFW5xP2R8dCWC9u4YlET2BXpebjPvS6CJjFoMpzBa0C1Ok14Ulqyf2kNX
v2G4K+33WTIQZoK1gjtgosX+sLz1oD+9TX5lvGGzkRDPeVNS53daLT0iACpUsd6Qwev3bBNVTTgJ
cct7Iyq0kYkkh4bAhBpiZSMlgcaCGdlhb5IJxPeY/liQSn3lnpqdB+CikwVWa35ihq4RMZxept4Y
AEXDXz9m/rz+mqRVUS2AxLPxCe4J7GPrYztWOj25uCYgAkiHoW2Clrb8VUsKwbNIxo3xBhpXdn2I
13nSYs0iCWzEc6QsGJN5iqrESrKPf3uMJldpM4t+6srO9906vK/xuwq3uVvOAqucS8X6mUBVINrW
mjHcJFyVRngTefKSmk9WwMkpCseNTiOPLpcSRNCutHDK/GpJpLmB9PTZaLYeW/11w6vx67nxtzgU
PTnCTfVmY2/6GoTz6MxD6tokDt+5lXHjxHrB5N7N+LHm40ckvDsE+iuFUPrlqmLtOVR1INYKPJKC
OjCYuTxtesd946H8P2yScWWq+0SmQ4SY6caImGTWzvO6sWOI2LGYvealR/D6FjKpry15PlBBq9Uy
IrPf9Peo6ZeQ+UyBjthwWOpHCOgiAJPXQjeEVrrxqZxgezsolAmQpyfw3BUZU/lpA/g/LWb91F3m
vWItlE+3icIcEFC0PuRlVv0AfK1hW7Z3h0ly4gusVDzBgeYJ6ggMsyO4REOYJK7+1YGgqSogwYMx
bwXGIil7aCW2XyST0XW5VntG23+UZTwqApsB+SIEX65VWSVzaNWR/nIqLf/OBAMtLSyWFV6cAbTb
fLJTLIFuN5OUVFDUoxR+fPLo9hGHb+0SDY0cR5wH3MUVdxOotDozbTeJ69XwWD6zpMTe+9xgkA6d
1VdqyGigDfZ0bU2F5eu6TSg32lHuUmVMwMSufDlVbHnIoF2ESH99/XL+F7rT3IawldMausfbDFU1
tPwy68X1JOxx5wN3xaYe3dF/ktLm0Kuslz+GK+sTvkJKp+CZ1AErL83o2GHjp69Olv/FetZrPjs9
RIAbGv7MqaKcuWmgLc6yF50vH/Mqpa4IW7+VgIK3jRSYbU0zZV6B0peKqg6q6yfdes4FlQRIusLI
UvkNHYohMNOv+or5R/Q/kDr7K3OXcZLVko5GECS435Z8LacbAkg62tMKDza8qROXpdXY+JAP45Qx
VtCtYVzl4bYcuH9J2ceJh/ttp6sWcPgOiwM00FpOIe0xhZczRMZNbhycPZicW+NgjiuGtY1HUAUD
E/hjQx7NChBET/n8dmSSeHt7+ce9RejWcZC1w5TqyQG1qXsFb2DWGsDTajpGz1WLDN14XSNVcQ3m
QnQJugR4e4tbQPUxKn1oGnnnVghhTKxNDkXglL9uab3cUUYkfpW2OoO76WHtJwvjbGQtlVG02MR3
U5KAJl6PzPvydgheP9uhc9QMj4u4WmlNqS34K7+fEscIKDGIgiEVwPuuEoEFCfMJGGDFvZiBTNAJ
l5nOAUsNQB75D64v5FU0R2KA9GrYheSyHkAvTsWIrF9i0q+p+bYXPgaZyqMiOhwVp5tsvsbfujcl
12fmncKKXAd/WGyqwLzuG/+LDQeha0UjpFdWTa5z3OfQWyq0bp1lyRGRIRw6j7v6TnhdnXYqPsDp
9Q5gAZ2JW45+73hXTDyphK+L4d0HGjiXfi1dUHDEhsSN6Se0xRsdqhOaz5WH8+uekeFWvne8r4gb
KUfFE9qlh5dW+yLTDl4rj4svkdsVLiCzQ+wSTscce2iQ4rQaNIEe0JbDm0Vz8vTpejHE1JiEuN84
NRH+BF4KV7MvcR8aQYA+L7odU0Oc79I5EaN5BDeKdMlNzGel/+67PVXbd8FoO6arHffzEcRfuZ7P
K6ye+LvaZJs8i2jP7TiqSAwFLVpeCac1NDmb3PalIMq4LagyMY/zOhcPGjwxLIVhT/K1lk4o1SBO
aBnQy66woBFx+CZ/070g49kSHhSCYgw8P25UCrX1gJTE0KQ7OXW/E32fBSfkNSo6esPfktKRbkbS
sGq0SctqPNwdYJ7hXl0s1Vy6urXAGwtC7KFIt5vLxP5wV6TB/ZF+PebaNZEGifkphg1DwxFyM3SM
kGSF3Fs9vakjSmyrpP43zODowoaCmhi/XcwJuPT4LTXnLPL6G1wiiwZjkNUh1XZJiKWQtv+C77P9
bk+rKISYXUCi4SITgQQRY/mjpS82GdBQnkOQOKu9KBkvuJZlc5GR0cBYy5oHk8RmAf0lLku7LR9b
FgrR+UMm1D0pgBCq3Dop1NGovFKoogaet97uJT5/DyBET9o8RoYUNBmJhRbFGNgR7HnPWWxz5Ch+
L7GnCdloLqjoODL82EVnQ5fWrNuxy5frPnzmdVuGEjbpSXD3ZYNqk/g/C12NlDYlqgIu29pAYVqt
golgeHFxbfGVerZ7Bnh6XZQ4fK93IWhRt8U+sfpX+DKJEZp1WDzRPUSPoVRHbTVDbvI3X0RBhYIk
IHZyl58Qe3D9iOVuHG0fBCY6BiC2ayVJs4X8vaxijMmpJ0DoNmgHdiUXBs77oF/9qWgnR6NaiTC7
i5NUXL/5R7O1P9+gjCZPCiewGJkUUbvnusUOuIKTNMJF0TOZN3QA750HmptbUBnYaCF9mC9OOqA5
7yqR/+H4DfYH45MJ+tf2eFhxMDJKIh1RgAqmnyTWs+v2mKCuRrwn2KVhGH3lf6zvqXaD5nnGM+Y1
SMbEfh8Nzwf4XGA6d7vsSRaHZ0f5A9qG5WKK2QdunKicBin9LtwNA+TITh7g6ahj4p1kNQ0j0dID
sOgY8JP4Vexg9GCuNLJiaWYr/XMPGvKZ4TPTOPzz5EnabhDllS4lkpT8JvxDQmxbnAqWFPGMKOyV
AcnuZjgqGv4jf69g1Lr/Y200RnZ4Pjl8/ABvm9L2gfacrY8GKQk68plXEfFqLVg4/wrGoVoeG6L5
BlTrgw4HFBOcSocZjXEgLNAhe1qVHOvJQqOCG7GX45vxxYSKvhUxgG2HP5YDcWNoYWEVLfCmDbrr
HfjeTtq6Tw7BES7GZCnsJ/CsFjqPgNc3koCxgAA37hnZGCBk75+hQRp2iyoUFw5BGe2leQrnpdu/
ZO6tMJWuK5HDz1Z7A6INf1K9TZQGnhUFkVWyRjUUrCVQmUEfGBFMcAd0h1B4K+N/RpksAjpGJV9e
DqividFn1QSdRphKbIAZL4n078S7TYVAYb6GvB9R6N+gKL/4oZZSE3Jm5a8FB3aXLR2HkZGHfMnH
E86p+Vj4gGESnyy6jFTAR9rF3T6Kq4B8u86pRBCTQ2E9L1Dnrc0vGoshI6zrV/GBjqBf6opYrQSA
StvbTAsVG6gveI/sWcnAJ1iteGa4kRYuVeHsaiMD23K6JbKGmjEitkRE+ytgEiojN0eB+5AyofBG
TPj5Fh1vC/nqjdKb177HsQSaFUgLAMTGaZ8hMirFxGZgk+CVLU/7oprqSefeEWcVTPzc6HoOXq0L
znxNyu+HicXOQ1EnxIU8DSssa2BA9tebmtfqTEvjvNeq75YmKQ/YRMinxCaOYOhMd806kMUWYRTA
PDrox/gNBbiRmzCPUnSgNorhb5SFZ5AtV/2nTKZbWRZMBgiRcKCl2kxtaxTmZeIuAvKexda1udN3
WpeDu1mS2/O6KWtzrTgKKQJjjjknJwW4KTKoHr5e9J5FRMUfuGJZjzSrT0VABswF+y2c2xz+aYe+
iqn6HavnH2KDmywwBXm7nueLJUrD96mF7iI/JzPoV5uDevic1ovpgzNmGobnibjdCu/03qcmiSBU
Bhk6mvAEhpKNfi4LNQyVcv0gTTn3agrxffi528lkAXbOF4I6zBI9hQOWlEXp8afNwfBAgMFeHmTx
t5g+5Hzfdsk7PjOWHj7rJyVOVA9Z/VkHUnIGszsP8CelLBMQX0jMJXELX5ej5Tji2AuvRQQ0V2dI
pvfhTMnEEF35qrwhEasnxHS566XgN4GXdHnHZWrSf5vqEQfLZIp4JG6EMTwDhXBEBt8/sBL187iT
YKrAzUsY6FiHanw+3lbtwFPGsecn1akMOviuhPh3VE4Qql2o5NPX2LEFg/id9KUlLvI0oRNkYe0L
QlVdNeKczeB8VnZYeSYUHKAZgi7Fc28WLi1Hzl7pK7ZfgQAIZEOO3tckTlqDufVnuE0fIfDjvDLr
Xtl+YQWpE1XSy4Qknw+szImAJXgZU3JvwJ4bXMzHwM53Ldd9bHQLugL/hR0z/5qNOn5ALoTzS2XP
NZllHaT5bcRaTcfs5zITaG5eAlV9F7HZnI5RaGtYUO61jATWKVtaAZ250BDYWCNybm4aaHwCVxXE
FG5+6VWsjwnestsH71UoodJUmc10ISNgPtePUwLZY6VfYhDFVLHkvbH3IGaKLh07vTQ8KKzQaVYe
A0aAoIc10KP0UXSvPPZkHZ8d0YD/QFeO/aqKMyLA9jtBDwMFPE9QMQHF99ne6HRYklN7xocBDUZM
fxYKjd086mltLhuerAOxCMe3R9N2DwFpj7gJZhqobRxv1nhrbD6OkYdKR4PxY8VnlnJiHK1CT12I
B0s8K3LdObe/676GZr2zxM4pHfKJBg0NykmgcxB9bgmf36uJDiGVKLWsD9aVCBAqSgeD0B61eRoa
TBy1REupG82Mhw/yiu0KMWiYWM4nI+WOR/f5jnDTrQsY7T5gmZm3U1XVUZ5PkgukhQim4miai+FT
ad8EAYWNT3cDz/L/XES0PYp9jr5lRqhA4LNFY6NMaNcGzgt4DJnFy/RVYXTqD9tQKIPnKvq5DPQV
yoxIzGGLXkVlP+vEJ1ZLpQJiRO0G3mvOXyr8gE9tNM7FGIoRcEVuV0rQ0S5AXN1mDNXpIe1q0+TF
b91G7f9pMdm2Ri2uN7kbeF2fkeg81e573yAxRZo6Xke0SUSleso0rLLK2dXFuoy2GvZ3ARxOMAOH
H3gFEEF/kL0RZuKUSzGmj9uLsJk+4sKvwF3cWvuxLnsuSUDH+Qq5M9H+FBz4Mb2krKNAj342wwSM
r7YuuVH1sjTl85oOtzlo57P/TUD7ADTsENOd70o3B1nKGiQcBg9tj1YCa6IMQ2yWvDltO+S0kbCR
IcoqfDu+Y6cs3fGr1iwFHA+Ewp1VUnGqlY69v8qMOXa/qpO4l761omF1P+voqzH9kn/1V5laTAtW
aXPdOAJmPQRAZlp7ZmstfzcGt3NFJgEJSpkW4CNncwGtMT7tcGatUtHdvGClw5JeUEXTyzsMMoJx
eIiido/I6d92MTPqbn8ABfheKZdCwHiKup26wWwZDvwg24leJVjAfXkqG85ZZGhYhO0wzKpW2Lol
IhkT6jmYsn9E53PSRa4NBwTmetu85K1mrQ2r5llZ4S2ApfBzA68nn6eyemaHJMz08RqkgMqWWL2I
HwEsi0TwClsqRin5JHYVUHLzFYFYi/aenfFE59leglcNeZfEE6l2mBgi0Q513/Zc9A8a/RlcYV7h
5p4SZ1sf6AXwb+kCJy/plj2pIethRa7NTF3vVGewKepMgRs/YrVAJYR47DC/nhX83yttGiMWijUo
qMCIQcIt+ZErgkVRQan6lFvSCuCi9ES9aXxnA7j/Xy/lq2qfdKwKUHdOHaFMvP3mizLvqXluqSN1
NIy3boGlp2f4CLlrJZFSBKw2Z6SULpXcCgpVUoasDPIyZVFcgWzrm1X72eA3GxAbxfLqrbgxCJ4G
v993Zio48UIc6240qN9gDbw9dNUj/UwJdHjd3lbsJou5lZyZlLIKzXncCymmOGqyxCQgouyqoaQK
EtKSVZQu/6FCUqswvZV0mByQn/pVsgBqYbAplAs3Y2A7Sx90QTEJbM+1J2X0J7f/3Nw99KgpuVvX
pCVSq4E+I6XXWTzVfgfIwOSDGKoyubixMDX+WB8xRIxPmsgkpNZ5yRaj/C6DYdyJqEnZETH0Xbgf
Rg6+W/2MHEdlj3V0v3nSZ0VKoXNINLONfEkuZ66KyPUY1pQegw594O93kbFz2OpllBb8xVkaR0Pm
8CVFvE/ePwfazIOkn9ZttE38G6eNlXcTrncv2r11MTnr9ZfUvygwfTzZIpEQ9Ya13OVVW3hgVa/1
RhrhvbDx9wOA4gO+1Z3d70qTHi2c5reVxR2E8jf4CExbquRtmzLt5mLVTgotbE3jlQuTiOjA7jxX
GC4aorGc1NrRHm9PwHnLR5ZVYj80fASOCO96p+VDN58vcE7c0kA09DqWAgWc7GrI9vLJLJE4vgy7
1l/HuguxdGZ+yFCwT5OsQcuKqKAORSz+8L0L9GvQGm+NVWwp6nFn6BV8DG+a3bebC9YrO9AP2t0t
rfgDx0Z1sK8lTsQBJv81kSGSB7BsKYK2Gfta3eCDbw3czs8DxLotr3SxlzHztM+YwCBJ4fdYOelA
Zo6fHe9DsSwTxDNX48Ej10ShyzPZ+oxaOx/DEj8z2lyaPff4Y3re7BRUK0slZrXATP1q18YGHRzH
Ua4vZHdVjIAvWhpeOAJhUjdKkBd6W3NZJQkiKPZq3aXK9tWRc40YRZF9RXkAl+Ir26Qk/HiIfsnW
/UchOQZP+7BmEn9P7DksjhP1HJxrzEC1r9YYciMyxlTrJ8/QgvbVgsMR0HhnqOlp8/RgfzgI0zPS
YqCiiLQeKWe25c21u9QzCNRt00EOQIc+9oN1dGbr7ZmqdAffptnVdqCL6Zo2Gic901L/58O4Sc21
deeN0tpe6BHm+FZhZrlUhzrjzWHdNvdL6RcXo4QUB//uVFyxZrgKW20dwhFozWr7FuS9Pm0lts5s
/pVStSsit9uhNFO0eAjFMh2QOKa/1FDVWi2cVT7jnaFliLjzKQBchIhgzXQW3Hpin0Yw7X+4RxO9
jokM/qD4hBBA+QVzLPsPP0Dw36yXzfRTlhsJdDKazCmkvWBRfrb3ZNNCW8PpMWKxtgMmrltncQto
jGxJORm846T/0I2/08p9KMpW13G9DgI7QY3G+2sex1bCJGuYlO0bt5Rt3DmRtyah8PyiS745Lmr+
ctHpSm6kmbBEPuXp/fkpqbrbP5Xw6ZERjdA+8GKjhBLVscALtqqIXsw2Od+768KN+LFiLToRVM/v
NN7xaXWuJRJEDjsObYmHTbgiLh4zcmxJvvFrreCcusgkyNKVDDRYimG/oqFtMEGLe90+FWR14bLG
jw8IBD/r/+U2kCd8Z2qm7ss8Z4KGx9UrcBIB8CAoOlpJUOGacOBFprJjX2p/4W/qka/MhzF7O3Ow
AjKN9FoTXsbQrx6EzN7IdbKWsgdf/pn66awhQzbA3c61av+Qx/wOL4x48QRvmxYOS9WsA6GKQcMc
eLflqSJfg82XtpsgRVMkCDmbpmYkoEeGxGegxRcXGWH5VgmDcDs6lTVNt4NVAOUNGJ18G63B1LkB
0lfDASrEJsmh7gBpMvVM2LNJbIq1OZztTRA/xnBXv0SjN4xlOzE3zcTFxUvxM/Cz14n7AKs1Xc+2
ZGvea7saNAc8zQBu8H0PKy+QkeFu8prUJbBX6GaDkWnReBsspSQs/5YK5v1P8KI8nKJdfswSwPjF
wyjE2SW8M2SyvbFvnXVV4hpru8Zy7YESMCSfOj1oB6uhJngpsPbjxjtWAyF2/11tgosnZK8V0ytZ
tuCTQpN19Q1gdcDX4vFBgx/cUJmOTwc9NGglue5dCb4yk7UIwFfABrfd6FWjUhbqHwDLuNd0rHMF
YRZMAa0/sC+/q3uPzFYNLneSbYsmOGKscoy4kI92qhhNfLajBwl/s5yr7tojQhZ1jSEe/pQNrSw3
2eItT/BJweQHeiG6uSXHZFkQhTYVqKYpcmbu6Pdt3L1D3x3Z9gaU2bYTRF1Ry91VpkvNHTLDHXcY
tCjkWrJOrzJsuGhqz4Vv9Rq9i128MA9mkCSWkHlb+xYbylpuiLXj+ccGW6pUXbatgUY307J9DUBN
Rn2HyMDCRwvQWgcdYZF28fRu1ELEB4fZa8deAI4YdcPB6LZtEppiJeGcG01NwxHwqkzn6BF31k1O
ypFCbLMtTJzCXNmAO+/2QDkE7ns+8vG4Z13HMrNzILVvV8voOt4OB6bT3jcWlZsIT/garOy2qxg8
DtH39nujc+ajQPvg9SWiDaXiC3WXD5AWz9BtHO4JeMXb7ZWpcdKpxRdqMe4WZrHXtA0l5kBPzt+8
U0tKYkGrWs+BxA71qQ6vHCP0UIaxCog2cdQ0nLekCUQ/uL6wiq/R+hAh30+qHBfR0aF4+tLTN+G4
sikXYMBofltQf8F00G2eOwloBg5/pEk40HLBTp0wG4o0FtSFg6wC2DDJhxbKhftyaQ4yBQl+q6HI
ntCnQvEnM2ro8TrE8ZA23XyA7EH/RFhfp0zNuLpf/A/Vr6Rt8vtiN2M3/O3e+C+G7ABczo8o3ziC
wHvfNPMyJIPX3+qcf7xS/rz5L+EuchyetvuFmKWR0BOicCwFCUYOo/trHLcpvVK3tz0vURlR9Q3G
p5IECSMkXtDyuqwNwImXD05TYGqI2CgJ5bAYCxIxUlZFatLES8RS5S0BMzCp4kLJ1WU/3WllBIaP
jX6Qf3/8Y8M09Do9rDj47Wz9zvlN4EkStjWfQyAF/+q6ouJW0Ok6xnmaMYCSt4OqwCOSenYfHN/Y
CFS6pOtrzzGvHA3pX/t6dvY8GyanBlQZAtn2NDn11uhX/iErfApa8E/NsEtsExMDM+6M6VjVT0gw
kauJ8cREWx9npHCFCDzPR25P105usMTA3TSJbEYbXRGOFKdo9HSb9mGBr5wolzm06QAPuYs0Hb0S
JXUcYteVoLnHtQ21ChOCKGEjuzDWpsb+r7fbO1BETOjpwq3L5aUUvR0oRc0PvYYuxwj+Sw+JRJJn
cVu+uKlzLB+ZzvfbEVJDKZkTcF2xGHnWLOMHQg1TIwq988hg7MWstRE2k6EadAisPKhXOOFURU6N
YyVGSgt/Jp/CwcMXbd8KZlFG3xxH+B+oqmxY5o3NaJRkU0CxMril74ptXSnYXEpb67/2G2ys/p/G
eEN04dYBnAVukQ0Hui6wt+RfLxgpTqXQFEOCJ7oUQWLIsuU7h5y6viyhtlBy+e+D7UsP2nv1Urvz
4AP8aAOmjNxLSxSbrtLSSEmmA32qrmYbnbQ8XonIFXf/dpw5cHRQxquSs1/UeS80Qqym1p4Qe4jT
47/hORBF/bJkHMFRQ0Qw2CANF6CemauZX+Z5KZkoDRgu8B3uhmRPCcCn2HLIDVdOJY8lRkDABNei
RZ2JTGx7oN9bPovYDvarolXPKVcy0lDJWXv2pTZDhd34AmRGZWjc9RP+Jo2jVwqwUT8qd6XS97i6
KQDKI4RD+qKcasFP5tOfp4TRe1Pp4FLJEkVWEN9S6eZYTzCrjRoy06HTv+w8qvL95kOGFt1E46uW
pRsG8zRwBYZr0I7AiagKf/CQ/wh05xgvU8jTnVAB313wfxK6UGXjBeMkvKf+BWquC2QC9B72Ghjw
P/fASTxaDtEOZ+AAOsPy9+lYFlammfFW4E++jRoDthzMCAGevGe6LFR5hTI+BgBcK2GiFpFjEOgp
R5pdEsp6Z8FmO8yRhr6hrZbN33cUblEd0pW6HnAZdJlPgOJlbpVSRH0tDG95YKrW8zNRWkk+d9cs
myUkuntAbI67lHL2fLcO59bkNq3cDZuU2sFgAuFlQecjROLfg5U78MiPqGDC+Uplh42tUMxRJgQa
1Bfao4AK7UibKtTqD5d5zO7CIFCQ63TdcMBVytVttkHzCOEGZnIOEZOSVonbtQohOnWfyt8iA5g1
FiRnFmSCBkeCo63oVIT/VRWa0/t9du6Wh3qORnua6ySjLswi/rP0TFoDdJlcSFDnLaJ19r8EMRv4
/N0MUkSqRdJfglQnYqjWm8vVmex74hCAiFvoUZZDpdTq9Q/rdfNBJZXtYG4YDS49TSYb7yGdrRjq
uC+NJaMZegi2EjVIrvezVE1L5dJwm7KTjSheuc/0OTsNthNttnFxXO8eusPEIh9n/nA8sWVFyBa4
eXfJA9eeHLUuAAxsbGK8KefOiPjRat2ABCc4XLTYr39tFItUwSBedeRkNCMPF7v7WW5BHGQ4PoOz
H6l8eviTz+JNXd2G+TuEQqADnplctMzx9mIxfUdfVP4+yP/DDklnrwOfyKMXFvlE7AUV9Qn5XsjQ
04WhVH8b/e0kqgDLGpIgYQTeK3WprysRa+w3trHpNdqlXdneJwyspop3Q7zSvLWaSHyOcBgtVQ0G
nGOmVC92bzXRJO4x55xYwF63C7TyNdsoPb5OgPjqDju/A2aeO05eJ7IkwxH2QyRECf0E26jgfQQr
EbCYnc2A8IzFtOlAu3lLvDiuTGtxZqMK0vnnyILGAVvOCVmSmSow/5Kw75C3SxsIXPbHLAc7zJAW
vULWcfJxTe9KDPjvwlIC5t9lz/F99wlORou4Vi6daeDbwwv6ZHM34reBo2jAnfiE+W6uqbEGWEGv
tkFC+wIRx1WwjIT7EsfSSEOsh9dSjrT/F8Y4bP+mmCA6DjN80aTHf9qUOGptAiNidRTFroaNC1UM
qzjNen4UjoVdCw+RynOyN5aN2AKJ0l0qG0tqJVKIOTy2g37rrzVY6fp3dQu59UzkgDyRd3nb+BL2
CzVU3HspAdOI1C6JsJUCuWtZ9pvpmjm3v9Vk4hyCivinkd18DjbPQ5cYSF1ZS3bsY26cSwyCKlL2
Y0IlhPUxLnoMhiO1rvchNZaMyodkJIrD/tes6ETwRUPrqHAtdArAW6RL7312k8azbm3ZiROdbAbL
WwOS6pH/GZhWwExcZt1mFTWZCaYIVUgduHyAYLKQdh0T1XhHsVIP5efHNKgaAw4rUPHlAun75Quf
uBOjbwKgOW5N5cjqwf4Tatzb+J8gTPVKnfZFt8Zl+dmfFNTIXMrL+jYgmV55jM+uq4wFVj/+uArr
qa1e0t0NjLEeXl2IzCJXQlulOXkbZZ4eqH5loONuKK4KGmh00MO7by/COeFLJapJudMSfJPKmkO7
G/2ZL3gNFcMc3IUc87b30Bl/VrZ76AnogqRacYedx4OwhMo14qR3RF7wjiZIFamgUE8c/yTjIfY2
KK/iuJKk3N3wZ4Wg7nJ1x5J2DGEMwjxtwjgqJzTDY4wz9IpdEQ6C8MMfKVtGITH6Bs+8MrnFYRYZ
AbfyyzEBmXzHHpTE+93XZVRInhtz9I42oe+EWNIHRvEZfiIhoOn5ekqAXSqh7TiEGw3Dp0sKfa1u
um699TmO4cA7drC51agsTHN05awWMup6hWlzczP98F2on4KG+nrmiDx7NoOfkDIdSpwNrBXq0Cet
d8tWB7CSxqObZb5962xOq1rgnOUfiCfn19g8vQNNjwRD1L0pArUt95ZfbxNuk5DtGR59Jhz6qeuV
PCkaF227Ff+NnamB9aZcU48SfDmy3/C5OvjG2CBnZIEjo3+/KxEiG/QQvLpc6GSQj/D3GZpjpZhg
Ag/m1hM/OtYPE3+MWjaqbAmWEmdg/V0CW5u2mQRgAbYwhh1+kxPsTCLrWniXJwBY0YNiE7h/fir4
pZ8LA52LpzeFSwvmO7Ov0YiPHd8NtsPPH/sC915hE3l5/C9NQMkGnrEp+18l/ie9/+Y4pOFCbD1d
K6HMzrWyC53N/lANe0pOpZqx1+LCT2IPw/AtNtaTs4hw0KejCZ3z+SbHZIisrVTDNmI/qGJxIrtL
7pxt+rVbyS/WuRULi8LgwiY8TP0K9EY6qzu7D0Avtq1IgifgNQE0pR1N5KC0NA3fxMxu7MWe1C9O
uJy98GbOGTfSrveX7Vwazuv4ZbFAsa4SRZQPeDDsuXuLWUZ9zmtwSquc5pkATmNoD3Qox/QpS58X
hjofTVQvu84CMakZ+hRl7NF8Aly0lCWCgGpYr/F/GzVgNm+5whce3KDgg4D+gw5J+EJVs7ZeGJWS
c7nPePxtTPLHLzGtPX0Rr5qt1IrEgadYpGDCsxw1jy/GNjNtKLXQ9K6uWxUj1i8bvMeLQC0znwpq
0VbsU4qZAGs4Hs3oi88fVW8WXufkgSC+gm3barCHA43ijiCm6+Wd9iLMD8Q9pmcbiPJawUr7aYRR
gMd/dMR70kF9sZ/Ysgo8lmR7SwwrFQWsgtOOrjKNuOKGR0FFPWiXvjlB0b9mXXfVQvxgwD3e0C0P
68EqDFFtEtq0xlbJJrKh/xg5NRLMQEMlw6nys6AryJ5oG1NDsITlsG9SEedKEnY933fUZf78ruTb
/Z4sGPMBjjgqHbQG4g9xvo3GiCZekv7Pao/+CEQ/tkXhO1FWCzC12VtKyjhEYmHVu9PW67RQKl1v
RyZYCf9uDniqzjNotUXz5GDJfqi0zKqfh7ZnMpfo//K2UjMaarQbLKssn1mV1jqHuesuH1qfU6NC
ONR/EGsj3oHJ86a3MPl6Ka5gFpyjXMMNU66i7MMBah8BJ4/VNsW/z158wTvh8LV0jStNOcCJSKW5
IDT+UExuV25MmPQU7rtoI81BRJY2ktw1AdmBrALsJSPeTCX96Kh5iJb6T3fcOXynoylKdAuGrG+m
u+jE8JSuzC/m/hM96CeXN/PnKeb3wHUaut2fK/0Sx06RpWfZcG3bxB2ztLXfQgv02xPwsAPdR8zA
u/1rJCmRovGKT8730nF+r7ncOvUhMLfblf38U5ZM+CPqDtwsRjNCg3ZU8AJQ8A8q1AuPL6ZTNQC7
bvq8k5RHTAeBn6pF47qTA3SBtUQR/VvERr+FnMi+nnxEQV6gcf5TCQRtVcpi/+rESa3q0wNmslR8
lW1ANo0GGN7YXbxnIdsclEvSaUaLJSxSaCYvLaq10P+nAHxUPvH2O+JVDNgzoVDKT/l9xWraJOBT
kUOUeKtKRc//46bIQtnrHqvmYB3zH+C0E8HHHTYGgoy+k/CZ5m8diZsLTcS2HXUBcTU0aBcAz7kT
ivHw4e5ifS1allkjUT9Zkco/LasNB0Ytduf5smEPJui9VSEXRDqMg4Uc4SNMe6+7puDmk0BN3d+U
GO/e9119+4bg3phrDBzPA+osjc6SzwHzIIdAVr6Au6+XOgnlZdiHCWbW7/YMU4zoANjXjI9h+Xwy
/hgP99pUs8S4Bc6RNKfrvNzvGFSNz4Uuyf2r+/D0+annaih8yHF3568V7ylo9hep0vVpuEbB+50D
g0hme3MysfNgDSASCyJ/9LdpkzklkIsC4Vd4USFp2HotPaDwwAfsCoeBm15EsFCtmBwU5lgU0DFk
zhER7PSMahpiCRK+a1cGXnwxVGz5Sbuz5WvT6yEDtoAJiaGtm58uXXn59gnUlw2/DgwSB3dAeSwi
e9qhMBmbJFMic/x8EcVdbqDEGnunPSkCNL7XOxjyCnsL6E/bmn39c/f5Fr3q+unCuE1qvvKUYF5H
ZHqotX/VHsxOy/c475r//g3wBHnfTU2S/ObMEorlHYMreulw+CvzgdvVrS8VZ3xe51/p0hj6Pp9V
cmBwVeGPgUhTlHriOVAJLF51VXEp3wQ3ScIoY5lshVmi/+VF6ZlRjB6qf1LQPTbeW4Ad0X1ApUfF
pwctIKYfmhnJefuj7Wt3o9ShJ03DGfkjhfNGEkg61/NogDiHI/AMBWCUpX5Od3B+LxCziNzVyRC9
4gRtGZfwhQINuVyv1zYAPAvx7SDu3T5nHtUbJCEOjwkAweYlIV7+8oqiZTe1cgsdV0C8QqQ3RdP4
mHYL2i+TLpW0yAct69i3nl7ElwxeRWfdIJotBl4RS2oGcUiKeVvvKU2D+ouc7SoA9+PcvIQG6tiC
tQCvnnejY/+1b6q9v3xr4R8XYMFhu0nbweVOn3no6GM7G+z1+b1TJRxHrSaZth3fyqBnr8NJb5KX
wbUUVHB5flN4Zzce/LAwD+qpsjlZ8zXFjrnD5OwDfNelfklkhgSw5cBVmBDl3dmZXjb3rW1peiF8
8eIh8EjoMjY/iqWxDp9CQAitP/RF6cHpKtzJVj1S/xLQSrxK7ZChIsXL/TR6IiTNLo+uyYibOzw3
Tx8Mh1OCbCk2rdYJzBOcUAReBH57sNx9u/VMIedQP2zX9aKE5AS2AhDgFCZwS9tO0PV+PXQVddPh
ibQ2UE+ArCNxj7cxCfEjVJEUkSahH+ab0Xtbi3XRbMDg6qS6DuLjsJ6/boDfulE6Swla6zy4bAKc
Q6/UsPXbhhTYrisKY3wtiPS5HZ8pScl7FnSfGOTHaYliinv+0Pyzsi6SyCqd3/lMI1IZDZIAeLUx
B2bCsbuYynCxxr1mN8NeDUhGo9PcwjGMBtIf8OumL+jmMZVvfXEr0SMWrsulwkRWrSn1GNfnm4u7
ehfYYoUiorEAvGkjTVP7b54LV2JlqFCSDyqFs/tUtMaDFUwkOVSyi6mXN37jQbaJxsn7QXxBjp0/
VNlNS0ruXr+ComRJt3W2J5Flt6+SuL1Q+otYnaurUWzY42a3nKjsaenoFyHzKOM0sGS+d8xh+xQW
KeCC9isBVP4WReXKR1hIaROiMGmxd3iGn4/RmN+8jQNYIPvfmowvAfeUkyT2m2w3ENonWKeK7Sjf
RDAmqNedvPV5djEA0EffdNPKE27iDZ45jOH1sptUUcVIQ9f14JxX3o+ZSyxCKh9rgMC4tkW9waXp
nI2ungT5dBbiTx4otcD9IS3F90iXRYX/8NJKF0STw5kNZgicjnStwFtZVNTaRI9U4yxvwrKAjb2x
aqTdQWm3pMsAAcscoVAfgSb8pYRV2QYED5uCE2UJHU9tL8zfgUlOcs2tGqxhdurVQido2Tl+nGGR
UqqJBFnRRT+288JyEG7Bew2o64xU5+skG0egaiSybTHiSxD8O/KTxZZQDdZoQwdkM5iPTd3pckXg
zs0qZq7Rlk5ezMZYLo9T1F8zFJ4HR8AvVzgiyuO0L7BWS8BDuW/8P3jgnB8lSMiWPnyS6zzZIDVU
MKBO+syZiAg/tq1UZBpEFiLMky6hx0JG07oUmei0QDqX4oEzstb9yvmlBRFHG8LsPFc6OreA8Ua4
NoiErwc+na4xTmjYGqttYfhKTfW2k5/Rt6TvNmlmSzBFkjtzwSNXeCIjdCZSHvLsbJKlQoRSLs9y
VQc7FlUuHWSpnxmrRR8N2A+SdU3KK85V8zSUVw5mfaY21J67Fk9JXVQhVZRm+cFAAZAlU5XJE5tt
9kX6szJ1bRz9LTfQPAUlnRuYDA3FP49KgfECG0ov2IXWc4Kw+KQo7sTKn6cfpQaoz4rcBt6H9m2c
ZISIWA10SClnJuVbqkpgTOKSZbATutO7j1q4Wnhk2BepPJZOq4EekkhrE5A5wvAFE/I0JQPoryYQ
7uiwj1QEmI7muSMWSklutlIrKrW9Fzw2HJ+yNOIMsxhxfSnlAxwzU0NSX4TcO2nsEOPSxaI96aMt
bT2YMpQXS8SMoicrZY8OyLCsnXXL9UWWVuts/esoKlaLPQn0Q8HdJsWTskmHq9v0hL6+jsA6qI1W
2bemjC5FhNpoFFn4A/v2i3Kj4M3rR9sthb93SVrfwM1040ZmOilnbFwm2cPSKN39gpwo4McXpNbT
0gmUM3Irwk7CkuoY5JNiygOxIZ4NxI4peD+1o6Wj0AtONSAOVAlM8TSsOH2knVnyiuYM5QJTXtHj
cXdSogSDhMgrp3wzATcZ0FrqS1du5IGQADO7EdF3+6mhi/mt2Pq5UaCL9mThiVAyL/OLPSq1V1R9
gSHKK6znLo/e78iaBQUpznzlQsTpvtG98LjgRY4zAZLM2q2zl9a/zM0b470vg5u1YTw73xdm5/o6
17J34ykojZsFPp8CzuepMdUddfkOnP3X6LwAZ6hHgTnurqlbqOsKwaJ/icxzbYremBwYX2j24HU7
tjLtCaRdkErCzaP3TaHYn3x1l3t4aRUjj2ni3LAhELW8XUa9bdUIlw2ZM7CxVM8QYlllvVXP69+k
oSbI1PVjT8fTCapW7Ivd0hAbhTtNORS7WqvTxuF8g22YxbxangoEh7EyLghS/VIxuG9ZyFF5a7LG
zALeL5WsC+oHg94OoM9SA6ED63Ab1udNgApC8YVF34yPZICEZF3EA9oMOe19tYHyf1Hjy4qpG+ed
dffM/uFk1LBEc8h241AE4zkpIgVOg7D2k+bVORFshOPozAgl2tUXyJnJxdo7JKdiEuxJvJOpb2WE
+qYWu82uIl38IOHbb1HmPxeu7/Fq8xBQ/0WV/xxaSBaMAv515rX8bHXrwkNEAZzn9UDpm9BIeDA2
9WUxLvKUvPoZYsWgCR2htyLHSObMy3ew28ferWC4qK4OgRPwMcpR0tWTkKTL4UqDfhoiKNQOfmzi
c/I2Gxd/ZeR2LcX+WdzuSa9OoXsUNHPwa5Vzz48ye13HFqMwFWAWGZNxWGGkpL1ViK4BX35jwwMb
WqcZuljgU7JaNDOpKcUgbOQoeqB7KjYPnAA6IZici9tENS/lqQvkC549CK2bwGWAXWATERKb6gMY
hVcN6+QErXUKl/mpoNv+G3Hwded8ZLcdnoZZi75Y9sRzb6Bqey77qEv5Xfnvxov8nWfgUg8Zq66V
1NW3LxlRvW/nO9lf1mVlvp/ZJC+AO7aW5XutWiqkAvQwXWbe1IzWtAaFsqj3gVewvgX1t8z8Rh+q
HFRopVJtxoK9wOWNb6K74bYTC/N4G427mapVGXUiYy5Sw/U4vUHKye/GjsAsytjriWe7QuLcaFIw
+y7cVD3pFM+ZEnc95o0p84IQ/dN0B3B7veU2GyeIxl+WhcUKLa/l3Z8T3xYBE0pZnvzFXAP+EVGw
+EpU7Zw2gJCNTLFWkDGvFYtFiQ7YOj5U5ZVFxhyKjyxpGi0rzlmnL04eu/6jfz/fAoPgmVCf/bL3
IAjAZ2e/+/VCnq2HKTpf6Bc4O57Yaz4QHVA6aBiocTYapg4CyCLp6s3nCqlT/eAfREMTGJ0/Ci7Y
yT/CH6WFYjrAiwb6NyRVB9NrnVpt/Vnzf+Q14z0z0NBAJCoYpFr3otASwVXujw8bKPVdjjIonZ0/
bdvAIl8OKdMGw18Kmm7mtrlkydKIEutoOE0VPEMkhkRqq75DjyEQ1Bw+SBuePEgu4dItCdflxtHt
zWCiuIqigNYb3jHv8AGGleDf1Oh1noJ363KvIA5ujSGkQrdGUTbmxdsxN4aPanGFCfrkN1SUgkfK
rozTH7nUy0V/JuYO8q8Voy3xDlgQkJsnZLuqhPiganq93qqOXkLWOjiw5bUPhqMnl+B2DRDyKPnm
lwNw3GCqrLCjgFsy5x6HIDGJ/j9ldW042IidQ9oNvoEZNpeAgF2z2Kk5+U7XWsKC/8pg5GNrMf2S
57f0nu/BtPewxaOhKo1zx5G1jgO1GSKCLg0yTACoVC9FBBsuNDcv9lrU+1MPLZ932Y5tFMNizARI
Oz18YmNyr45kMxj9qeUGs37E8zB1lqPzxS0oAM71LypNcWaK1uRgNLsetUrRY6+ItO8pHW9RvVRr
bF4E2loLEGeD9unWIMwxdohrg4gNrsOtRTrm+wfjtbUobAGKDQbuGNT41Y+qbZ6vpc8D3Z8O3+S9
kfxHpOiQtNVJW+91K9axk0+7p2uwFrtqfw+o8y0WHmveFS3AOONeP+LNT+R0oma8hucqAmM+XPd/
JFgy/K4+4H/fkJwhfa4E7sY5Ey2VqNLsf1SdNyJxMBdbGgx4/ki5v+vFr2vfDDTC3LFyWOXnnvgy
BCdkUPMhgB8WMnPinY8IjlAFvuaw+wh20WEagfx9sFSW4PNwavTHO6/s1M2vXsW1O2ID7UMrxNoM
YsNKF+DALKDhXHjUwX/jyyjEo4oNIsXWrDA9KEJGObbB9ByXW0GhLdYviPaa7+rSi19Yf59GmQgD
Uy/EzQIPhbARrhDUtZxObJb0brvhdHwM6vynUOpYy9tKBW779PUmL8IRuvtSsOMLYUb8oAaMtGRC
hoGWfRCg7QVJH9lePDmYCEYS9+5/PxeDAfnetltl4B0yyiYN3PnQ2vto8i0Qnj5tABNyeXlh8sUZ
GPDhIxMMYz9VB6Hg3KRXP8VyDU1ChupnXdbeWckKMOh2YRP+o3gSJKxEeKofVu7WPvXgMkYWq0l1
bzHv5//JMWBLg1OLf7hmI68OtTgrxDxwNpWzTZ3nLbEaLDkRL9wxS7TBzu+lxDT0V+KRkbeQpIO/
o3U9Am9wy5OcrrOwh1iGZQLR6/TrpVNc9UU+kWqtRTIxWQ/Ap7uxlk5NbtmhMwrDO0/I21rNBDUG
O7Rry1C74vuv6tL2teCKAeAXtAwessmcwMozenC7nfw41QMS9nNG5WmkS5dHyQCqWeRypJhOEAF3
p6Lo/3GZjqdtw/q8NeUPA9/APNepa60BunUK0G6nJBYTX1zL/SKSGIYYnmWXYBSrCpw1e3SEvf4g
llCfvgwEu1Nmwu8qPwnl/Tu0iPILvAayHxnsDJ7abHxvCY4rCp0uegO435lmr9zqykt3Mt3/s3Dj
MDwEn4KUlj5lJeROe7skZEKoXvrj94kAS4cpYgfXb22GPt8aJ/he90A6mdFTcOvBhNmRIT92jKva
+NtMfM3VqQyJpxuVZ5ZpZE5/qQL9KY2woLd9mUAedwE4JCOC29libm2nv7gp8NL+P3HncEAirPmA
WbeCto2aYmRolPxZdEfg37qe0+YJPZwL6DQDcJE0WTH6tQ+g1/qc41KPfWLJ2RUf02ojLdItR3+6
O2gZhYkpmr+IARknDQ+a50svrYPOjmNbhn59qwxinB6kDXmy4MCUmJc6HWCHAqfuS0MHIXN0A3IK
OpuVCCpdZWL06P38wYmHMgAjo32ypmaqy9Q75O8xNoN8DAF0393nSR/6XPDBjrpLEi8I81Xnfwrs
kEe0ccs0758Zb7EOz1Gr5vR9PowiqXgKNAk4PfW35l4zNpRZfEGi9pil2ZharhA9CdCElBEAATq1
xaXf57VMfIaJyNqL16twUyJ6U5l/UPLc0P4HNNip8e+aQWR9rXC1066AojSnqi2ge+iV2Y57AF6+
E87LMMp/BaeyQUopSnFnkF1Pf5D8EaQb9xiDWMkQPKDgFOpyV6lHXvDrVQ8HKqwW0XPTj9PpXOcU
3tH6K+HeDt/4n+g7+g/jg/pwS6+a1qS0lCGatBl1h9TvP5bj3Qq4Xma1khYkRkJNVnQ2bOHbEvAQ
oLQqd/naeWwuRQ5jW3QVBLEKMB4ZBuHRQ3EQzm9sahiMKE279sYnAyC0/rfMrLQhgcdo7m9Y/KDa
+wt8RQVZ2LjJ7JbI8dxyGX1RT/BnJABi9jQ2PXOTXair8HDMRF1mX+iH8qGc5kJSSHM69coJBzPA
3xjo9Aj1NlL38vagoQDkh85Qz9ElfsfNQlKh0z6KhCoFnAJ40WxBle+NRKyhYCBqC1cRs2Hd6imI
0PVrpukvv1tl9UFv1W90bjiSse8VhG16q/lW7oweSArfB6vFy/sHpeD4Ac0e3tsonpoPK3SnJqTw
0aaEgyXA/Fa8Yo6ShEu4Htl55Z1GRW1UvMQ77jS4PoiRxI3nyDtjnmxEH7dI8nfTQjVzBIHng9ZJ
ZZy2g4WMUXTbu2676l8MXYaydmrK57mlMM6PeIZ0xTRud+BiqB4Uqvuwv1LJAy8Rp3AAzAWDd3Fi
pxxOnRp82AaCmo6tBmUsu3YK82AzybRQn/mI7s7SekTpFMrkqT/446+3rfMzFNstejqycdjgMru3
4+LaWtGo/fRzfwvgRP8GzdwxyUxKHbmjrCJBZfe3sVUtFZbDlhaPZIUpEVaeS1VYb4D1Ak9n/DBw
UkhQuxoBrxtwLQOvhbyOdk/kJuS+SLoH3fvq+dsrD4CY7OL03k1RChmIo4UB8gU67QeIHoowBQNK
gxmQXwMq7HDrZc1rQqLfB84jSYfDpOUQfTDFTfk6tlmEwe2Owo8OVdHD1rBX5GVXyk31/RZ9g/TU
V64ZO3rWiJQ7t6AezgVgw0OqgvApVs8eRQeNk7SKhq/bg5HJ7qDZsBQ/zZpV01GNywbsFf/UWn4n
IfwoBWKrWhIw2/h9DmXMLfdHbokevKUnhTVBy7zkmruJX38eHPeVEUTQTUVx5+WVlomDX+QvJWmz
y+wTOE+U9zUlNPYcX7rriM4SCA5exuqeCVBsG3rQFoxlcoQTuqyg9vTyIas147Le2ldTYbvJPGMO
XYj9gf9+lOXtgwqoqhhMwp7VUpE/7VC6dz4ys2mPOeMWeprKYgCKypZVoDbQmY1W1q2gKhhyIGFt
DHkAUkVfabTrlhkXc1sH2eOw16f72dTGt/XCPdG0l/BtrwouKKH1WDA9PJlkrKq1aIXqkQSwgX64
r7ExF6bEvOWwfzBROVqaGnShxGhWw58rLFckPdHNv9x6t/IVG6637z+zC3+wSAHre7Xg4TeQOpIx
YCravtPo/SmWwlHYBAAMZaJl6Egqyelws9MtZ5+8P1sLhRu9leihnKdtvnZ4b78p3VLzsI2hL6Ur
+Wm1F9chZSkwCceSjhqjvUdmZEVK4We8bxFdeD7tfwWT6zcOFaFfgxFW+r7QtwD6UXpVNggHiWiV
DAHgHzTAnDmXQXtn5I07G482YDrpVZCR5FpprWm0UWouJm7zuYO8WnNYBrkvyv0Gbknuq/UTYnK9
xFwQc3b5jCe613zTMZA0pBVo6ynVdPmzJiyWb21vPyN9VFDCTqw4pLkcW+iADeejJkKG3/CkJ/nI
4UkTwEzpesWacnJ2QGmX3D3hrWl/ruMTx9p//vNZm5WxvCaXjAH3G0hdYW1VTBCZPgjRpPoGZf/r
1YkHs5j4u55spDIkpc+kCMdffmu6o41LX0vpSby5asoucYYThv4XDDifn+KB9bPWALVcueyd9UpH
960XFa43XVQEKWjcVHOfACk1qqrZXx8Dib22YE5+8MC0PymCI1Eho+U69SBMVVAXc4FPqpv1bahM
9canweB6XA/07DsUjBU/nkDY0Y8we1dW6ZS66FvV4j7w3/XTTKT9XTkkwdlFGjsYDVQkCnndouYT
2nMPxM/zgXh2y9CqUe8EROwFEg2/cGE8pMMtgTbm9mIQml39fWtyUqzzfInEIbKlz4DtCQCgifX3
jJuCGjyHsrGrKNZU4cpwXoheFxlvj3Gx02FJJlAfKMlfYZoxISVcIDevVNAzjZ18voTWCup5t/xL
Ui3qMvso/d9aptabAscrXsfR6qJnDWTT9YIxhwsBsUeQNK7ApDHw/usAebVRwtyuEUHU9LwaenSl
JEDQw/d/1EoT0rFV7n/TWMbsKAFWN45rFxUvEZdqCE7Bf7dHZRjsZgCSU12ium/7mGaTfqLAtASm
1rXYCU5KGRPovidDaHRQpOKbWULqMu9Oedvqeyu0b0lLEee+xtI7OP1TY1HcJjGCHnHmumt2BtjC
ny9EXI31fpoX+UHYSb3NY/oOG4F5KINZ66L0FPDKXbB65O/ajVZm7hrYXoJV7ndcE8O1PmUnYaa8
k8/3y3Bm/PYjBaBaa7KPMStDeuu/+7AkDmV6Ft6EV3L+kKu4t7KIVKHwb61gfpKQ/y2BifNF+7EK
CZGIPpBBqKPx4/WLrqZTQTet3Pc2YRU53wrQhdX+bGynVpHPTHLna+GjH3oxWsqcc7WGDMX5hkst
fZvXC0m1V/Tp8BXKys3exh4l77p994GXVns22ZwcvZdOU53+kFdyLh3P5FSW7q3nrHBCC6UMzuhJ
t9zQGReslxctC739mdoMlJhY+0qZ4EYW7qkyW8XV3IH5U5uknULi//IO/SCBPZ/ujLj68QTgajYt
uDp1W06ehrP26v66otdUuJzkr2hXs6MkioxOWH7mVxpGLLYNhCoktsVtOxGyeCeyxXrcFToscEyX
v9i7XRU5OyRziSJHDn+fyQiJTMFVk8UXXsroCsBzvm2ot5V+cw9umjjqq+8J2m85lH70irylLou1
d84bMuR1X3vPpG2Wljc+92z+iRnPgGBOKcYAc20pjWeY2bhm+z8NkGd2/tfHfsbx55PHbnPm908z
6c8IPD06u92CUjW2C6LZVa50VpO9LTVU/CDaJH8oyRpGi+u71SvVBuxQWioOhR+0h4vjqDcrhROe
YFAirzlG6suvCyplzR0qyjo29gHSZsrNcENGM5z5viHiamo2ZnTD1STn0xGdTpiwfpI0Tb2wZLOB
XWJzysZ7eZYoCgK79zkU2wowAY9KwKo/m0m2/29Zd7oMxmbBvZK0Drvno8NMBcKY+gnoxZnAAH+B
s7vESklt8iPvOnU0wMinwPHzXBvH90CNutMnwNxsCnXG/1WruvhMhi/IFIgg31z3wLgL2m/iRH36
qVcSf9YSGNgpdj0QD8/vQrvMCPv/NjVoypN5xnR6m8s6Otbyd0Yag5CkaaiMUaCgGIG/DN0G2t40
+fsE9dOK9FXVA8lK/mbl2nRq039ECO3w6LzCwImmgEV9XWIMuCXcgDfKrpiePAk3Xm61mx4RPEEl
eteGP5EwL1IFUUESQYGO7WXLTHVw4sN3RLSSTDsNA4wnb8rH2J77dWPdrVukGSIeZ8UpezublL94
k8nmgYOuFvQtsbbR1zECScEwpeTv9R/TiZaiIhuHdwNTTmcVY1dKX6Asojw3FXCoeOlLgYD0jO6+
oupmJns/GBQFnbAliEzFd5ykkLnWJTeEbduAzc05TEMc6A3kDvlrxS7yDcKIz+8p2eXlhduvgq7r
YfypmvVSTIn+lei+Nj8dGqnqO3vf/SdxQKnw5RTw1bHYRtYHyHFNZv1a83p3B6F939l/8FzrLppR
4BbDgsGJGaCcFy07lDG1NFommn5WAQtgTelWwPrAmfJ8AvOFejTdoyCRIBmV5EmUh6Jg+Dp3Oxij
f3JLamkSi9jq3yokZo2ZA4bW4SsOYRNuVLuXZb1FyNX0rhzBBVHhbSOy2bnEjz4nIRhNfzJtBJM5
CKIaJpe7ZkpwZt5Pl7AZ1TDhJ9GVCSkqM5yzhgKq/73Wh3CTkonDMhNquTpxaVg1hLv2KZaGEwOM
sIvYpCuUdrJ6017QtXdd93c6BK3iQXjDi+PNd4zY2B36QJ6/ebdTUYOT34LuwjERU2ZDfKfL8v7a
kCXtX7R/2Fsx1FTbDsbhYDct+5oT5Bd4MI9wO/I9oVkbivz5/Sj8yk/LbStoXOTFoET6rXsWxmPz
sd9lyAyZz0+siRRK/9gzcdW2u3lLMmLds2v9l0SGNlWbNajn1n85+tmRgoKo8d6Cz7pj9klu8/T9
lfkKVv1sNPJQry9Y0pAogW++FkZmJEknZA8WqEZlSF9x1CeSlXkNhWtfPSc+7sCW8rVXYZNJrlhi
BGw+IIFXxfbHkeOnkMNi44ip74+uHhIqHkuD/npWpX5P3YKUYvbZfs+fg+v+AeIfxVpYJobT2lcG
8VQUGBijqFYAOMZ05JaemGXWjIPctuX5P3J5pOy28XcfuZouSazVG3d6O41eVde4/cdfaSNlil7K
GjCNcsdpbdo2NUtPQZRDEPJAhibNL0niryuQKRHAqsk2oGJV0A86I5EpF9C56lUgykhXzzvA1c53
J3m/f9dq9OaRtU2dACSF+f3qOi1lCAPt8gWpyLzFFC+LrEDqC2QJYFt2cLGmJ6Fx/sVFY/hfsnvj
RdLN26b9dDUfe6jQDHrhLaAmT6/2/XJ6puo2xDaXy26pz1AFY/07+fegcBhA/nW3uY48oPoLysEm
/dKVKK1NUzw9cK6WwibD/I2AGc5VXnHqH4SvN1X8XPNu6aHLKlRybcDC6nZnrUCeeGdipJc2j2Rp
FfHcM93eNQtEo0D1ew1kY3GQdOnd2P6r4Lo114HEv1i7N3+bo2HzPTy/i19j7m7h1rornkzQ2NRU
axpQxQcdn5teLB8XwwL0PgJSa9NVpUkDBBU2qJt/Iy9QcaPssprBWnSjQNJ3OyEriZ0MeYOU7iFz
9RQRtpEJhE71/1I6dUMODQcrJsM1PkpAng1FKx7ikahJ4I6PRdlY4YuOsD+sftX1j9l3rSj5bnHZ
QMXGmlBqFM6FeZI9RqgLGlizQu5ok4m8HLhcWl+fNusnk44E3RJPlru8DfB3EbhmdEWMaXs95PKC
CPtm7WWhgsPGykwaj8f7qC5UYDyximSCZJJJLYnMQmUeGzOxMomrzznjNkNGeBwN3BcCUVmq6PO6
0XhWcvWUrm13LkFSw36YnK35Plaoa3O92WaGm0fCHYuXJlnp51tt8ttCy04ssP7uRfrQe6+HOq4q
u27JBpJ11QseyDkt/GQrbdILFqGXZRHMSUhYAw8XO2ruPMUy1BjkNNwcIKYotvp0nk3PU27g00Ey
kXm5Or6J5xjqjw5lovq+kyHS/Ejoniace1fkEVTZ6kTfC5+KCUldEablSBuKyqmtaNydl2URLSym
zcofn0vCU+Ip+zwaXUlZtmIfaiIoMsYgFFKoFwsxe/roO1Hse2SyNpGJTPtmjdoIXAfKR3+goTKg
4hGf1UQ7swVPdGNhIioxlNDdobUNeU7Xi4eve059VSjW0OX7DKrOG3mJ7Wzxx4Xwt6O1xIAeOsEE
4atmXpqMbUO9QOVeRcNh7m5wgw7wlPKqA+L4YX6yYDAP7i0ixbFQynB1Ccla3hkOVDu4+ZKN/t9T
Zh24aqi7j//RaxWEIiQdI4yWOcXiRnCDRLBFREMc0vo7aAWl61dN8HCsS5A1f3pTuuQbs6ur0vTZ
T38ny13/7LJ7xJEPcNqZwU+mWy/SrqPSMRAAysd6ExDiGyGLsO6pHz5nje3otF1ptSPImZ7SPyZI
3nyL2lnaXvWq1L+qf/1Hfn+yJl24pMdhOlMULiq5Fm1D1XWHKw+Q3pDl3QewXvqxFtbqDVau9nZW
kd7QHa0ENtV8ahfggQXotjNmvOFv1A7jmSbZgQfJDGQGe3JX3zjYRHHz898y2Qc+RD/8rM+c1EMg
6xugZsJ2JPl+vJuw0CAjgMmMlcrsc8s/mjYTKA0PcW7PeQVy6jsQNs7RRbHeQD2EfrcsZq4GY07L
t7eUvLtBpXUQ2Se0qj5DXea8Svjn8lC12vAwDQnrX24iOoZKlgb/8jM1014GzJHHHeVHApFWEWpV
SlaQxOhqPyB0j5t8LiUk3ig4uCCgmzvEMmGAAj2v+Tco0XMCoxki0J5DXMRbVQ/KTr321N/hq5jN
ejl1zfdcW1c7OvYMAEizCiHXW/BaInH7FO65XLO448BKk2kyOE31DwkBBNK//sWvnRbxmkFEt7m+
0HVDPsZDnYyBrj4nBlBMlYz6HdNiJsGK3pa+HwXbF+KcdtqlwoDhIMntP09Ydlp2E0lsCTGwQRVP
dejbQA7SorKGVXl0nr6FSFQi7vwmH9eSa4yd+kJSbs2YlpmniM+9roj31j1qfjmj4AUkqo5mxs36
6vkeCcR09npm9QPs8wGbicKm7GxUBRhPIzBMUPVxwXs2XiwAUUYtGJivrENcQarlzbNiDOCXPY3n
5odtlRoSLYz5OiUQUwNFiWRNDSDEQFHUjht+O/ZZrM1Hp8M5XZfhNLA2udeVRsjT5EPcnuKoMB1j
K0ZgHEM4GGSYb0B7hKhdxosChiF79tTBAUGL6JAGPFG/g44n6ip/lrzl7bP5bxrAZxdUbkH0BfdR
sA9lxtlkUCkixP4juPVBAcn1odUWrS91PfB8IrIHLZwML2UGVr2+54CdIHU20xtyZy+qbgsJritW
GzfemdLuzbYfT9/yEz/hJTOTJ1gJqHowF2n28KdCur1ADPqXsHrhoustRu9E64Edew6NQTuZIdu5
mXT9tTryKWI4o6RP+4jp0Djh8UCA3hrnNPRD1pA+mGFSyqkvSzD74R9vLgf1/DNrHzRK9frusgIo
0nBP4ZlxKuIYYZ8mF8KZjU3LULfu22Xpv+AKFFclUM7hBcskbsL7TmeveD2YP3xiBrQW7fy3EJXH
x7e6vt+Rc9jhiX8cKG+BvmX4fOcJ3dm0+WS1bD4wUV/KhpBVA659Ekfo97UFy27Hn8+QqAhGzSiv
wJiUjigEblcvspiajw1UOYnMB01TR0s1OeAvxhtsMdeqojnMnftfX01xzaTMWvS7LUWLYD/tjTA9
Sc0YVup3IbRj6We/LxW4u2Uh1t188FNk9jVgV4eiPcXOhaR7mXCyVSwTD1LmRaNz0+T4fpbMPdfB
CkxMEbS5cFQJHdk/nwFqn5XpNWRjbKSc9Ly5/VYwuaCFLiU7G1KuWtozdyXYDyN2mNmEnFAeYthI
OvLxo5LNDKvaFxBR0bFuG11MnluOcKsYlm+/0jtsy+gWsKMUwwwiaW9LGHMnz4pjCbVnulA0q/bR
OJ6hBOc/IIQEA/2L3q+I/Kd71t0QGNMJiiGbt/4BDcngvKUh4ZlvhK0p8dBVmvjGngjg3eaEiX6Q
+Bur7eoUfDh7uzAtm++jqmN3Vw/md/t+5F2d+obpYJ7IETSoPZazfTzzbwuFbc2YA2lU7DPyt6br
v3sz0srdEPPRLbvDRRs6ODumr7SrQxvfG0YFTPJh4sNYdoO/PAJpNAWXPI5hnbNPY17vzgKCr5Nn
PGJVm82+4oDorWvjbQFqi5ayKlPvmwHSKHem3WBiEhb9WS4cRPQeUx/qdLos9ZL4pzia7kkwI8Fg
QDBgiQlMXuFif2lU3HLmfFn1Yh3yKge6EAMVnjand/Zt4C3DKurnD3ceetTggU1MGXoLniZ3s7Ef
n/0R9plW7p9RiWAEmKX+h2ThQXwK3mByHYZCZY1v8agKTzay9sfmliMK8W1RX8h6LkUo/HLWSIUN
/hdqmNz6AN5LJBOw8NSX/Fw+PdkyYvC4QKzO0xhi9yITd01ERHCTZfVKBsHScj2iZUdLx0CFsTRz
AqDyF7i3jEopbsWE0Y13+rXQtgrlvFJabT/YeBlnS0UL/jA5v9VXTfkp70J/+KpkgH95tdobFvhE
BCnNXZdyUYaYC9MPntR09Dte4bzuTmxD/4SijQbE0mo69yuxys3zfRwfg24VNfyqYpO5cXx+nrAT
Esi9IiVs5Zadkd7VHzWtkqXPBL6E9w3Qn8Ittvv/avWXfcW3hCXUGx1PONvtnFfc5YQN54W1qpoE
UaWeDQKogehgyikzyFBLS5309KZmh3IfvkrUfHhcw5u7nTzI9GKIEwV40/M3rTyJtkFM3TnUH/gm
0kSRXfSVdcL6JSUY6sROPvSg1QCrY+QhxfEC0uJJKqNCoiQahQEFRpezEd/LQNNspQq2fKrUkBgk
EEHCPnkTs9Qna4qE+Fw//zbSmF1m9uydOwL1q82JYeteFgZQ/YXPjSMI5fTcCIXsf7udvMDv1r0H
c52bJ4otuQ4hTGW9GrST2neDhrb02IZwFJRtlbkEwd80uek92N3L3g55V9nkKjyoCK9YPaRd8HnT
3x7ghwiksXucLiZNHxe83aHI0OWZKXo74Y8PPI9MJ04FeiA5T/j0isSGilJhoqEyuCmUQDoQVq9T
/pvjKSGRtELhR/Pj9vEyxt4rDXMMGT1MJLJ3pMPXAj+yAqjwoMq4kR5Htzdv31sXbQJoql62kPQp
Edzz8fFS7/IOTu6k6d7pRoKy51Z+CSnzwZt328idhdNu5qOpkgwk+wlTPwYI1W5pWOdXmv+DBxud
uYGAA3WZDNXDwS18YfO8rOXK+yY95XG+crvqR5ioa5LXShbg/GaRMm8iNT2ctXNHWypDhfYTHMGB
eUXXqO9d6Zf5AVjZNpS7WRcNnZ5nc3ZEHN9djVKSd2eBCgVF0LXF09GVES/PDFoRD53f6/wkkVIt
vf0K3v3iRM2xNh2JP/zKg9YeCvaBVcaCFAyXn1ySI3NQAwnhCzjXsGiKTJkhdm5YOvmm5XNrjKaT
IGnWr53971b2FPxSYVu2/Woz0Trr0eFoAfT5beoukljQhk20zgQqd3VWD0djfWLlUlfgkySZ6zyW
Xg0lf6qRD6hItXQmG10bYpjvIFkIcZkQwJKeNniNSTZgPMaSLf+5JjZ4e7TfI8L9GprW+UBsncul
apWhKOLutMFm2TGk72iy3hZJCXjA/QJ5Sc3LEQZLjcAZSuyLiG8HZVg670bCyxQYwn3r6U9XLN5M
O9it4ZsjUgdS3FchWhA5bjuYxgOr6EnPbBRGwUbVlNF2nQW4l3cBZliOeUbhaDwPb4SrUWL6csUt
xezeDmaWZhldlo9LZtaMJdCqEcRYESenk/IwQ56ld475YUjtkg1KDwhxK5O5EJJHtXvyrezNIkcO
fsmRGmtRdN4k6RgVD+dFDVf+qsI4tjAhIyEYSiRD5Z8cCcGETv2b3xaADs22g9ZfPMX5vL5fU/WJ
PeSjXYCuLkFlC2TeIs62lXCExllTVZTnLRNJgnGWNJY8RfNZmieykw8xUsdAr/wzDPKQc2jFAnrV
hoWq6USrul267jMC6uLMCZ7WVpW1YDUsFPz5Slo9TflQrm/s06a3hnPPKVhz65yR6C3Ucb3NFcug
lpnOs3uEbxFH9sDE9E9pSKCqNGcKpEUdc1g6o5W/eo0vmt8tn5Z4lOl5r6XgIGU+p7hluKM1UIFk
AsUpEE8Lr/KFPilJnnsOF/wmzSyu5u0clzULSnb6zg0BtRT0NA2edyxYNlui+QDeYa8W9ThAPmv/
v700BH4dKqJoNwxn3gSuRig3oQd3YPX3ULW185V1P44/D4avFR2uFphzxy8yg6hLv4VQhiFjls+2
wRUf1ziD1uAsPEnVaHTX+FeQA5uDCjvUgpIx2UtAIwSstws2qcBQI/awIdLr0Mnxb8ltR7v5iDo9
bDk9tshpx9aUC/xdckfK7cPGUFouLTs39ZsDXX5/QNTq5T8XhuHHdeuIWCpaLF/6COxC/wL7+A87
qYuTkqjlTbstV379YuNDRJDJrl3bAIWpi7ypSMMShWA13KZitQVnrqMpeAcRzl+5qiye3ZXqjJQY
okI+LrnYJqGFXoTcVHowO+Z303lnQR/CKIDXMoylI9D0Di30n+YupZUXEQ5b5NUA+4qhqosl9qjF
4V34eYkwTdBqp5IpXoCqlzNhXS6pojv9F7c+GwArh7Zq6K9QxsPPkbD2XSMZllYdnB1NJq2gPBNC
YRq6oLpnoBjq5lJwtxmRMLYeMMXCKbL1iR7+8sFZ+0SoOgwE1j6vhcjDGrRoPf4H69vS3SUOJGZ6
jcDKaC39nAtV+maNp8IjN219Kz9yTk0cb5PRE5rKH0fid9Emtavkl6hurUmcfxW5MJIvqrBq1BaV
zAs047SKuCsyRx4n1TXoWfPRT251KxL7XK55hNq9VFkd+t4vrOjdaM/QtMkMMcSQrLdNRoHKxJIA
bw9LMBHNP5zRleU/wiTQP/uRnk4HIBxwqLZ7dHke+ekyvUuiWqaB0k4rZ/6DCZNs7VrMUz49/gZ2
MPYeg5ZgjEQhP7XCmIangd4AJlJw+8gAH7Y5KpZoo8DcHal8R9rC0wAObiLpk+OgpDiz7y5MoB/l
dl2FzlrGe2djBVUmvQPyGo5xv2ns2xyFZXoQc6wl64CO+/IbvgU/r4jKO3tsm2wIYVvurx1Ok5A4
mMUyQ+EpHR6P+4eC1iA1KS8BEKSIqLUdggYvmygThMFFaejl87m3JZI8e/I2qqd27d/jvauNtC6s
9WGkgGpS0its8ntXroy2dKv831ysO/xB8/ijXUVeYrQ2xoyXAxwK2eNgyy5DdlBZ+kMqftK2lscp
Y9F1t/UjK9XNoDSCHzPQlcmANTO1pZoybeVVGBjtGTm8V95IGN3YLr6VbDc96TUXh8C8M5TcU+zq
SGNaVUMG3x/ZhlFGV5EtQRlF9DVPwgIVII7+xWYzjVgtQc8wTiNT0gopCRVoz+LCc+N5liuFaGei
DXkfGZp4XRpNlBZuTShA0X2MQNc/X5RCesZL7z5ehNzIB0mrGjGlL58BJA3hu5rEHsoZE6AxwM7k
tG7jTlhc96W+oovCmnTPNBd/phylxBfhMOHGhwXS60vHHpsjeqrgE+YPT4cd9ZM2lK9bkaD+aATw
MjmT4/2LrNLydS1c/A5ALcu9fUCYCzhqebpSBHB8e6UKXJYYwRNeDSJs+wieOhEGeveA0JOVzhtU
/AchlUWzkWRw52kGmpQ3xgPdZYbmc123MJ+J/otPWxQ6B4PnqIkEIDF15BhP0z3tjk3rBT8xSr7J
rOcoGnme126q4DattN6e6b/DW3T9yFfskkli6m1dH8pjk73iQehjkgG1HFLTOSYZawguoKpOJjjb
5ABtnZX6WLpDY/zt/c2SeCPOHHP75wpgVOSPLdgsPSxbsbzO967g/dgorgYhJd1dkeJl25k3LNq/
hhM2SK3W0Swz/VmKziGxHO8bhQPrI1kCAltRstSq0wwD+EpsMOz8CUXft6d34puJcQ0Tsu9pcBor
2Sjn+jtbwL57thpjOA9EntULCcG4GWCkQ0o/AFoNrYskKozE4ZWLqJE/ipcvlX6qL7CkVzbcmBOS
s7Y1O/3KQXkuyTjtTzfZm41IDIS9ssis6zP/CRXOoz+wqGp9D10AknIj3dIcY+X5Lr+uQlsn2pSt
kRijay2aXhOC4TDjTFnBXaNP4O6GuDDppICCOtkTZDPx0bZbrjBY2B63SxGlIRxiYVNyjKcfaV+9
Imw2HYGLCghxDMOP1Crwq1PPqTAX4UHq7YsfNYfmMBo/U3sKRoVhMxmL+ppG4XxhJJdZMcfVcm6R
X+OmzP/284rgu0Darw/us9nd3MqJknAxVGLvWAJS4ROzcPIaGDQQf/A22GGnRBvKevkvrj+XTucY
pxzVlYbG80bVi/nKSmHOrn4PFiFPRUUsdImj8seyv5IANOeo7WLCu35BBpN4lcSdI6BhRxJA4xpK
2gZ6eXJD5genJfGfJiNLekRUSwsDrp0GqTh5CKiGYIULiQci2QADIvzVzjbLbIbxOONkoZ/PDnRM
yCi9HxGxgE4O/jvuqcMwiF3HY3dFl2MhiW80v6K5x2bxEINf72RvdZw98HI13UDTkyHQWhRmqiZy
G4+BFQB8GvpYzaYtAi0s+uQzjqgbU4+8x/rCuyP0CSEIcUVMMXAX8unDLvO55oUnOgTNBkOuxbZu
jDqZnHZRhC1abLe6Derf1ZOx7wCs2ehAXwV3qbem1w1H5BsjlSjYlr/Qgr1dUYnn3Qk+jct9mVQ6
fW8iWrDtLtsik0xo1CDYaiHj5tWdHx9cWKeJ/SQAxZbVSg2SOLRvLBEsf7XM4HznIH9gd6xeM8Wh
itynsbDezkvnX3q6xai3GHelWa0TDk3ZBAa7PPjJRlYr/R+kiMKSYshXUnlSeIaVftW8oHgRoz2n
AKWtUAGLEa7X5Hf3AupzrdJt6JipRcDIW+yMX1wWh9pnXVvZHGJj1KGBVTYtUzXq5KZZnntfv54y
KOYGtCUARdAFkJUmr7x7j45wQTXVyvwl2qNepMhgoNq6IrQjGYDXfOg6LvUYVHvjn4TtWaxSV/M0
LYOf29lpr+IPyWa8QhXsnt6LiB5YCl5JyrCH3U3irvLxpEkKSPY0FJi0DvoDSLgVWaLkgtIWGO2L
H2gPh7LEfCb3MpnoMUCmTfev5Yq9SAvh5riavfSMY5iTFmrcUF33AJ9GFIK5p/9e6RLMXNHv8M1b
wIezySBfEcY3OZD69bDwuU6n0/wxU0TaarA5u9FYJrrZWkZbIIIkq8nOdRyL3NhZlnGGtYzBG60o
LlRZ7qHPt3AFwfOEm7T25i+aGNF01bgpjmcfI+TYIU1vNzFRF7Ww9jGPyNXI7v71N9PfugxQv9Ci
0i+mfkx30mkFfvlE7z53hzbJamUZOZEohAG5ChG/u3cz9YnIcGDz5GKLDk2IfqiZdI0yFn8MjTAL
YOq6zuV6RJvl+k8mFYmxoGs8YDvCSD06EQJMHnvL8PfbqPukt3DryEMHfqScNnif2VFm9NQ70C57
jnkkKhKAOKYgRLSnNfl5X+Lsd6camJg6PUEljxfUJk+NyJR7FNr9cPNpuZxIsWGCOMKzRonMXWpu
rVyEV5FA7M94sYsiCIb39Jzofwo4vAIQDSp61jpqucFG4xm2eQ+MfYmtCkINocacBVAmaWTw3cdg
3th2Oc5ShUQ2Eo8sZP6/T9UMh4S9Gg9K50C0cK7u6N9tMuoWtOU3ZOPiuTbsuO6dDGauI6uXYlyj
XTZbBuHnLr9SRIr4rO1s0OID9vdvH/sv04/ZD6vxJgF/K0KCnadZEt9DWlZtwphJHlaHBkCpmxVc
erQI5d9Uf1cBrDjNDqfXTnoFyD+zjSTtQVla/QBgahevGaqPC2xZzZ3Kc9MUH1cgb1CpmcDvlovm
MnOrXNrAnIX9CuaIS7Z/7d8b3RrALk2JuPOPtyIV+VNoL32931LFFVvwmSV66xU4svLADMqBwjSN
FBG1TTxh2QMXe7E0X5Tf3RcQSifZZMGFaUU50qPKwfk9vi2OeMKQT6jWbistlu5RouORUQ74+uxT
4/+SHvxoIQNkyDeKL3R3dAJceVntJV6lGfc00QZjS4Wq8h9J2ZlVShHq3ho/32nl9cq1OR22swtG
JpKban4T3IRYRgaF6Ae6+GIO7P4rwOskuoEMmdDrFAANtnpZwkm5IUulk3xRpKHc3WjblGjGP6Kw
26+pOw6k5fPrA42XkHY2bAOgoYEUJl6WIpv3lLEHalgXF1ezisR6KcQ9FQ7xHP+LedAN6BZZjtzL
pbk/h4uopWtZRqcdmUKsAewe+WPu14wZUAZuY5MFxgz28ZCXjURqHFVwS3lqj0uk5bFGXg6BbQmR
247dSXK0siN3WFRCJlnWnygbdtZ35LTClWYveuvh1mjI7LGLkqmV8xt4J7SsEbnPizkW1OkK7JW+
BP9++P+EYRKuzoeAJ9/GZUTQxhhOf8bdnzLu8Sl2k7F+gUP9ukExbD1pN5oN85zEaditIYeZQ7vr
ajUaCnZ6F2PIT/IHWqI7Brq2sHG/GCagVrCL33eBCanW3ZttYO26x3RfgZ8lFIuBuC+a/bQcTCcx
mpJZOLOdRbDUZ3f69lNrfax51cHXrU19Q0VjgyMuJk3+lyNnvjWKNP5nsKrmPV6o8/YkiFCQqORj
1GaFwqj4VeBnuJmAoobgucxJPx6mRLxDjsOmc2YdQwLoDoGNihOrJpGf4CW4oMWjtCuBTiqpN/jT
+tsoD0JrN3Nv+r2QVjEWgSnR9TlUt6gveDdKBfo62vGCwNSGsTkXGYd8gadhPlegYVC2o30426EV
D2QNsZqEya318R0dIgJeXwCty8lID9dlekhpnAoVRgHXaYUz8AU82Fwn37ABeVNpPvswmEmaI+Fr
9LYy/LKlVqyQi9Hgqf5gA/2voDGRRRlQxihpXvHJJ34wev+5USRQdIBY82EqBD4tdnRUpV2/TtxO
28fHoaO23mE/9BUMvc04yeFWuMn2ZIQMymIH6bf2bG16BGc2YvURS9RyGCnB/64E/VAKO6MUgSMS
jd2bT0V23dNtEwinLnFSh8ob20p7ePFOjrSjiPmCY1Gw7TuaQN7cEg/Jsq7XZjpRyv8ZkZAL8Uqp
uhTu1xTEFa3FrCLVb9xHYKjD41T5r626AFTq8sX9AdvH4r8te0TXjwynt51nKfwr4NxpdJi+rM6E
Uyo7EqB21O110dvDV2X3TQza+s2LYsu1fTDMr+p+OU2CrqvryMyQA+b69K+HEYqf53BE+MOdeiay
kGqQNDeLGLHrkrQ4TqahAjjxSixbA/JI9l4ofGJQVeUh3ezQKOJeL+e7KEDyTwraTmN86UVjaF1U
NBcvis9DjaGiavUZ2ww4U4Qoud92LrzUZVQqcCvWSEGOTk5atTUI9TfAt3pDTwNgDY64BnFWTVdI
91YxT+qNd9x4zneoSZsaiXm9ueH+9X+zn5fh+E2Ax2K17t5yA5FW9eJ5PodVQ5n/GfiQkBDlExzt
SGiYRvaH5OjBml2BGabC+AP7K8cIZyeLl3p0eGp/Dc8BpXljFlQbWzhIz3PPKsMRMYI0jTK1tyFi
AQGW40PS60nv3d+Efq/pYZpMjsNR9psfaLxz2exX1uf5RhVDdaUucZFsepvZJCdkPTHlppqscAZZ
Dc4249JPuz1yRK5qk8NiGTWOgH/WG0GTQ38JHB5wyDer24SHlCe6dkBnZzR3OMNiKT/7HjTeoK1r
RGzhP94DlatCmKr5xiO5h3WMNTT/IdYQwgyvuQ/OuF7/qiAV8QqTJPNBqstXkkEKgM7iWmDhnz8L
L0c/oEzrFwuIvUi2lLGahiqg1xITa4MnmUFpMLV6iA+bvKhFD2PTFKHA3tS3OKcHTvDBsY0IepQ5
4jPmvgIwA83yuSbXBAJjhpRdrD33If644FDgh3omaMrDqaQjUSvn0evY2SISSuh841iglkRkSjme
WYMFN+q3hrnhAwGfJnYBTCAn1oaR6YFnjlGiRt3NfKjYNLs+G8uPKQaDX9AMp5AAu18SlRdE/qjW
kg4qZ5ORkfStDRC676sg253sH2nIAmqLcM+baOr36fdCq436Sy10V8vlBgOfOpIXyEeeFNNoewHs
gmaYX2BUzxZJoZEan5Qr8HsZaQXlRh8LoRYc/sKZKqcjIOR1V4r/otQJ+p/VoZX5S5EqWLnIH3ue
Gn1szgousdUKGFS3NKTfa/9/kXIR2iMsZ2Okb6jSERlq/lnLCxDt2C6m7mPqZXAsqJzsatqjb8wF
+jkbYvChqTahJPQxFwSIYIauTsz+L/GgaEV0nyBdmxw4ReR64suaPllfUrhucfgK0r5f+N17jrlx
iuFCx/Os6R0NN5IL6YdeoIPSb5Wk1QUzmF6WQ0V0he/F1ZXqMK/O3AWb1HMhP03V6M7/4hT7HB1j
knDP8fJZhB+5H6TuOXYWulGjsHLoVzjgshFpVIbgqAILme/VxEed5Jb4gEkGC48WjIc53UVSGaq9
IcXlqb915NhRU6/kZmBNFhCso3nu4WJR3Zjly90vE2rjljX0/FxK6AeqfKxK3Rl16T4wCTHluM3Y
22+BkhLma6e7pk1VwZk4uvtiSWSFdfi3NCgogZ9N4fH8uRSeJH8FeDJOyofr5WQD2AGjLORdsrTp
5BxRAqcbcbv4Qr4T1ezs7CHBDSokef8MA2x2Wshulp6BvEVYLHl7KI2PiVKqwIdjg24Kek+O4xHw
/ja3PPUh4Pwn3ZExjq+hE1bxh52kcC2ls0UA/BF/GP80XChIafeKEeSjUVHdodi2HHSZPBzLcO/B
sxRFz36JhLMqaAZFm4eHqhs2bjbNvOksTCnWe0lsjQuSTeDFUvha11iPVu7R14x2Zr99U7t7ctIG
s8+74tNvZmfPl7OGkRhFGWhX0ZQvVDOIfFRPXAcQUjKa80wcjNIgZKqTX+al44MKxvIeBuMNWyYk
PNsju91tCOmbKNAK0giJD6rrXw05v1d+6eyIBW/TLTs2NUrDR/FA/l4mWyhOJ5y+JtjdyLMsnzUp
9y6QH2Xcs7J2Xu7ubO/rNDhqPG4nrkTi+J9BWbKqT/r2kUAv69h2EB88vYuQTC6noayxZbAxb68+
FD8lUgyTikaHPHYypngDVdIo+khMFEP4SBaN1BJO/KKOeeG8C0qMxWN0z4uj7+KsrbOGY+5yQ0A7
zHCxX96ayflp1Ma5aseAPncKXaNutK50gbRjyUt1Gi4HDg34WvL5wR4Yvu2uvT1GC5N6zh7TYD4j
Qlv5AZ0GFGhTqrfhhIbyohgfu/9gWEu5yPTCYFaqNK6MqhNd4HnGELLVu0U+yuuEghw6+elOiMSK
i+324/KYCEVDEMkBoDMZUgvmjcfUPh1gNnUenhPpWT28Qs7YBpcA98XL/hoqekJWVpe0bDK5UiFj
20kdbNbDeT834zgdkmyRfeTdkM0jFNlEmWSlAZNyMF05ZeNKA7J/CydAaaf0vAgy0Pif45AxQBqP
yZtfDKsm40/sRrsEszhHO3VGIG+nSept2fK0bhDf5OmPGHNfpfSkzRGOfUQwKkHVDYbyfmI2WYMO
BFbg5nIZSMN3/VZa6FUnADTpF/4/yz5Ig8fjeP6HM+DUJeeDIy8iyg+0AVJrVb//+XvPO3kou6Qa
p+tnVmU3/t8lCFS7ttnvbH11yyktWMe9v7j6ps+PZ/JughPxlhiA11bBN196YmuFg0UDTfuvDGEV
UJ6mSvgc4OQFpHnI7gFfkdT1C61hu9de2BzALjNpI0Fu8qdMlcrSDBKw+P7rC8j4vOtGxYy0hIq9
I3wstFBnd2DPINC8y3a7z4AJ6VvcpLn9F22cfDOaQYE9WcMSx9PeMrYwUT189SBdccKsuIc8iJl4
fm5CH/sbE4PtDBcsZ5ko96ZZ9FVrqctRCEFcEv3zOA5DiJENXg1Q1c5e+IUS80N+Ttb0WOpB4Usc
GOuRnI3vPJU/10c9CfIhiWFXlbch0gWfMzMXc6YwEuvnZc/h0zFMyIhlpP/kq9QVDkBrT7cn+9KS
Jkj9Gpf8ymZVxS6oV3pPme1iivrRTpq8IhM/MRCkN0Wbon0HJDuc3b88VFkc+XOIv+iuz+O1nYiS
uS/VrIqPyLDcirVF186zndsntkw8cqvinttZiIhPbguSzS8NV2wsLBzCoqDus+dxnuSJDLRJ3x2j
F+vkkSBViXh4bvWuxA57a8MRy5I7RlXatmIdstm1ZEXmgBWovHe7npl5msrRmI9Y+q8Kv9tRpw/J
A2pAqgmc/0V8xJ1h4JBK/uTev+M18L0yo0d2o44DVECoanSLCIDPqlXDZMRh4Fk7peD5Sw5as7am
FD3kGMZ3Y4RmEjvTPz67Tm6utDLTPrX9Odxb7oLisWpWLnMJij3c81zWaMyJ7/kWzb85xwa9sa1Y
E/Wk5tCl4I1tbLIlujQ4JHnPki3Dt4uSd2LUMkb3M5MzP11LpAIdC1QcofQiSxbgdZFIGi40IcL3
AcvFboE36bBVFaYh9HABdwQMRg8YcaR+bgMrcZzfV2BXaA/PZ7Z9WV/cX7ul/IdXITQEl9GyP8+O
PRtXoO8q2T6Zr2Z15xqX1bTG8FETU7p3JwfPOMLGi5ljFsTtgxkOKblQDd4Xo+CSdV3+hmAFt9JC
xUSKu82IqnYNosAumAb3l0KmWWtb2pJNESe6mq7AWpaWO7rk9HXm4wWN74jcHaYr8xPQBItkmkMA
yQPojWV5qxU+6jYG41Y151QN6QuDue+DGW5M+A9r01/Bc18sp8157MeA+j+zBfNxmo9owT0THWvn
5sER1YqfO0PV5LVcf8OQ+hXS1qmTWqnLAPEqRpTfec54v+Py1B43PFA+GKSsajaexB68voxRQVl8
8EAiGTvGYFdWv4l1eBoLRoFlL3Z4hKoGvep+9800ek8x39WK2ckGamO5DMWKn8ceMWPvu8XGVLTP
Mp3e6ooQQnBwUiloqYVCxwTnfharCA1lCP8oIAKfqUv4odtc8nqAFR5yW+8FrIwb/4SWdgUUH0xZ
EM0ychjDFMtLFsjvO3QfbFxyUWtIc2ryQxOlnRlUMcMxQ9DCJN5/zVLjJqwTbDGLHZ9gvMHWT5P3
W7nAfHRhwe7Y7sXmdAgKgAtKN8MwSv0/XV2bBUd2bEpo5jNoCwcTbMhHrstv2T8LPrsdjmDwywEj
RW3kokTDpbN9O6FysSy2YZ7HZKr5QSzjhUMV1ZQ6a/d7rpRCG4uV3KunvXyuiH5lWkX+H6WUrNsS
Nwz0imQOKnvRWu8/N+78e4AHK0AVUG8+toHVDFUFSpGlrlF0u7iWOxu75YKtMT8vaNba0J00mCS2
IfYvz5G4ItXPyEur177W7TqdMhaMfS2StufzRlAKYZJppF0GHvLcEObbhb6SynMDHkueZ8XBASIO
Cp2LIMpH2v0+Nvh/6JQM3gCupLHsspM2FeLV049KydXNruyaDyBrTMwZPpai2uDMMKNvjL3oqHmQ
0VuPNmPtdhRJY1rlJLdqJp58KxCogYhNwUfHpaDQlyWgwg/XL9A/fq4984t/MEXTzJJkGNachMeP
ELmXJFbpDJbEut0eJlNTflu29SJKdtCvyPfYTBSqwQJh3YZaoB2PUsofAZ8loebY/DUvIIBifkdS
fqXhUU6OPfQk0XFH0h6BI+xxyFAm6cmAS/wxARcE/UPRc4t7PLT4YORTKMf6njaGDbAY33rraZD7
60ACBPuEVDxjJRz+oExwPQOy5+FlstWiGiKp9DJwf65lFkGfVVOXxp91RaptVWzFVa1WeDc0oMNj
ggV3qURe9Y2JD3MGLSGe/cFLZwz6HeqzzeaXI3fFxLDBjqtrnbEMmCyb/9XCOwjdyWL6eQ71yHVQ
wo0Fz4lstjmx4C+PtP+p/wqWOnqE7DAGCYWftxkZrP4uKsK1sn2hrGnvyBv+oxKXbEX1i8mMM8e6
uhsDVRU/byL0vZJE5iXvUHNbxuPtBPCMoHi7yPZ18FYSL6IBBILNDERTmTBztFHOC30dsJLkSCtr
pjDxH+Tp8LQzhp+ckREl7NpsgnRMMPMgfAXNipfWEo5r1rC0h/qyxXd96GSpOJrCx9jjKDXGhrOB
/ksApVhjo4Il4Szz88EILQSPbWSNQcGazBJvEurRuZZvTwefCWkmjZoIAcuBVZjjOS5L9qd5jNEa
6i8fEF8vbmoH6h1P++wsnWxxou4xQtx8igRIJDw9NiaDROBl4c7Wl7PVEqm0lL01BQmyBqNHWhy2
A2cGdGKMxAFfXN2gAlSNhjLlpMCYKibEa0MJ9YC+WBpEeN8JrOJxT3PvC8dbNnkJoiPDoi70cc0H
aw7PRw9QPivSZKteMhBRVCQSJivA2rIoX2WhIoeO2SbQmPj8IboCHSIzXFhzPD0p4A/yqqh9iTq7
qXA2S375E9gISM8g//Yug2HwU4wK3ClV48p9vX8+G/vY9ApAeky7NdeJ5gcROCux6gCQeUxJK0WH
bp++w+Ww8cNLLex+T207woJZK+P87KNOj47zcIP3jGq1fk3EA7ObVboZ0g8QoSb5rpL2IQuUfohC
uKOSWhO6TqN24CRTU4sCrN6AtJi7PfX8aiHjS0zxP9zvlMfNocbK3lsIHV9B0YYvBk3KRGSQhFZT
Kki/2CfyQAaYAfk2dFISl2DyiwOK6EFyxaZmV6BtkfpfnOQ7zUmppAmalgLWMnRplH3sJUUtSWXa
mSEcWrLxMWrH8Ja4DMmKyM+Sx3QFp43szw8IVtFQiKR4QqmPX28NJjofroIELyWmueDAbSmqwm8G
5zAf6KpWSi/FiZQ3oTo3sg3QEe+FASDdo05PHWkdUxJ7F55mEjDv2BrwerbIXJ3oAEtFoN8Hh528
E4CHp/v3Tmcd+xsdIXxWlzBDyg9/lPxlb82zHpzS5GBgudh6tJEmUKcO1yF82BLLG25wX2y1thGd
6KpRFVgq7eGg53TzbUKxPvhiaS7OfsQ9D7lUxcw+og0Xf0NHV2TcT+bnNOw9meDFGLYA2tUudIvt
M1njRxjxL5SO+nG5UkCIu0bba6VIv0prGjaYsXDlP5jLcxHk1LYjMOO8bvZvNeVTBWN8OEIcEkNQ
aZm4eePhCEvBWlS1+2xdrFWN+gI0viX8Fw8CkCprNrx2nPWsVO0KqhXv5tYndX1Kb+l3x9fi7Tih
UfQKqHRkauA0FOmFEKjH8yT44YPEGPrqI/Z/s8r8JaWOZKxUg2/F9jmRcUintK/tu9HJtQMpcG1s
9oAXs9Gl6q+TKc0nUSzVB8QNF7u0JyG3hbXHTMMZ9qM2trjIysBZ3PY4GmOOhAelsK9nNqtrKG6P
U8mjBzT6JHUstvzg2pnmAOEzMwWF10hTfVeAUDYQLkX6p2vDRWjS+biX8iTTUVesJhO0pIRlXc0s
ABpalC+XxUh/Wn4tmV/WmnjHBL+FsSt5u41V/gqmD+oBQnP87o9EOk8yATddK7DPevQxNWdduFu9
kvs3cj+23sGj3xyemFy6QrhBSt36TcU6pGIaqk4y3zxNg9E7id/9Nu+e3befNJA/haxMBUZ39Q5A
aolrarPrTE3oAkmlYFiCj5Xvxpl1RrNMCQv859c9XprWJpgX1kNxapZz8PJQq8cQGSgOSc3oFGtc
ZaOmxSGpKWsmM8kXhW+wBBEB0/8+ScykmrcIeScVSlO2AbcRhyjUo5sIlCCKU4V4Em1OEtayb6SS
idhakj81euz59BIzfkvG0IXVsgRMpTRuaGI92Wsz9HZfc39Zrt6qV54iqM6O8pOUigbvMHv+95dI
UXeYfKEWTLeWFnA/XzoT8lFnkXPm7qNROxmBFb0tyMAVAU73yjtIyfy1+7IBwIbf3UkrvPKLwzJu
LSJokGcuXymTzgr5/wcq63b3iTzvNbSunJTa091VtZld0mKMzXeMeYavexMqXvJGY4Qvl3LCwJbC
5Br/oDXaSdvbg2KV/kjOsEq82Ntzhr3urYBPw9wTbwtGprlfE5lz7cBSVy0rnRKPs9N9w6WD7RKr
VhmWcnDWeUglWQ58hLrjFpX1ru6SQoq2CfW+ryA4xKCMl5wHiWU6/BxVF6PbQ4y/pcIGjssjS/y0
49oV787OYQBHlhfacVHIct0XKWSp2IuoMHSybFzlgXMfXatGW/ReeqIV3S+OrQ0+O8DTx+Nhl98+
Nv4zws7MC5Jk22WnvcK+RfoZZjI5GRDM0+44IROfg17K2qawkqeGKv9xfMZOQCzrF4DNRFQaT71b
NaUMd3pAGgPDpWq07arwWXWi45RpgQbTrXdITNYzV9JLpb8v4I5fODvjGC05Y++JsxS2g+3+c5nJ
WhHGFOsvDouNoWmLGXxvdl2wuaxhCfe+7DyOe83SfPUkbBOfffzvlQ3YPomASun/Kvb93fiu0Bsh
0Jw+sHehGrnDnIAQdc/36s2Z6zvN91wLKvAhkefH8qu4kGrp7NpoKHLTNb/8IRlhDbRCIFm04C0G
nDZrd6VRnryEZzxPHyXKriKDEGswFp3RUzSkHQtCRNlJVAZn/fOa/+xpmUWzVJ2QGZcLkSthrtsi
YqY8TnQUhwE0VVgHJsHHMI+yGlVOGBTTfSKAea4aD2f4XnSvtiZTKA+qZXe8DzPrW1eggXjFpBnK
rAJCmTEsp8SLLgSNjKZCltQwWf8kL7f5NCpLU8hxglJ64JW0FK+JfvZkNL1S/e3FAKGRdqOkodDn
Gwd2nQiltssGfXxE3DnlyQiYIpX7Zg+cm/STALon9IEW27KbHSQ0TIHrfNEUP3TmNT8mdPSXU0/g
1v/eaYi76AbcGs/be4G2pkRdWovA6Khy804PvUTUsS7GMgaGrsUTkBSQWNJSU20NbFYtuDMhtkUc
pAZ02iDkL+onSqRx7jFPgJmrSyoX+fzG/6u+Prwoo3NiAAwESCDF4i1957ZJUYkwCqV67mfdOH/Q
Ggl+01z3pU2+vlrut3WHPT4F+q0x3qvvSjMCx71wlXuKgbP+XM1aPGaE/dYHvVadx5PXeRHaLLxF
RRzgzyFRcLaswMcqYWv1ZDPaIWunmlwDKFFLkByJM9FxYPfCv+ZcHADj9+rlMWCni3b6injGa2oN
uoKNOexy54MFuJpNgcsojOzpxZKwUNagmog80wSLPvDeSGH/dqpUB83NEV/Qst8zlKCvcW5x2zrG
CqN8lZbTIHoH5u8HbV3SbLljRKAz5sHx0NPHn469JtSXR/k3L5nzsRUgb77oCnXa13m40IrFk11J
PqKSl9YPqgGBviza4lY0/gIEMLpXPtBNforiX9S1H5Thu2TCQq5Is+4NXBhHkWqED/r4xdZoDw2g
MsdPgf/UB7avw8iZkuiRGPYXG2b1dPTHtK1B7uEtKUdIHsFl2czJfW0kuDRH92joPPsT76USyfoa
cg9DzLLj3FrduGn+2XF/AbkEY+ORmDC/94EcBaqBAoue0auDW/um3en12/H+WJQrlwNhpVrLIBHb
w0eo6KWsTo751Cew9hd3CUkpxiD+NUvoSui9JJrzYT7gAdsBUOQf83zPyKSILdWZSncoTuypCsNQ
hxZoYsrnwL9B4g0ry203etYaO13++yf5lIHUK5Xl8oOcv/qnEp/xSDEjcHNxLJVKRqXPZLizYm6T
xXyN6cEHKJSJzr+VU6GbkwALYvXRoZx9j/G3zPlpLJfcQX5M6DB7Gei7gedko0PaTz54bW+vCPyn
A7DbSkKMQf1EDeBdzamKYGCnu1Hbiva8U9gU7BwUgAr9udbV+ClzLsZ/zYdga8bo3uUpkLR2vxaa
MC4aU5APxO9YdOu3QjGoLzRVwdTGoJwyti8q9G9J57sWdoygqs7Pz0sQfJcdQKXwFpQpMjfA9M3c
Df71m4g/wnjYDNcrr61n6d2BXYPRp/ot33dUrkKaZMWEfOFlZL3g2h1vcEzPpuxirIk+ReaVWkVL
BFK0DfjwaspWYkctzX9EFHHYtAmM8ayIDH2xMGSJLYqVQXDs50btrmfjAI6ad40sYJnT+bulBaKs
wmEAjTB8KbRUH7+WClKWngl6IRiz4L/qDUx0uzSDy2PPlac3qz4Re9hRPcGN4VWM/B1YFLcc7UTd
Y2mIqludxBgmJyjIfSwzGhJK7j475Fb8JU4qVVeJOqda2PGoQnMpg2YrMERan3kXBfiC5k/9iiKU
AKE3EcD9s4LqgoCATIz7juES98z4n0j/FGuuR+Otsa+nec5z/OWeM+zrgzGqjLP94Dr9qebSAsi0
CGnzbCuSnORkp21Y9bazJWBLvYFixrNxiwQYw6A+SaEH06Dw/YgkzU7IzsYTInACV7ubHG3VGzKE
FHJdkT4lU2I2fAufjrMmdwgUdqQvi/csn1SKB+fCX2V0nZhzpkBG6nRrXmZHLJO6eFcgF9XqmcgW
kcna6IYKx9fzabtBRlHRl+6CSi+wnX07mA7xEnOiIWm4amaElKjlO5SaTAcA9Aa404uG+eNMSf7P
t/DPJ999OL9CjX28255cYoywZPjE4M/JnqrpAKV28IxUMVnuzV2gBlAUA8Z7jL+NvV3yJ+8hnueO
4oZQsvpLEW7zErDEIlpCswZXQO22ORvKKS44h2neqx7+LNp5Q7GHoBxA2R3kFfUnTRb0Id2mOB6G
bpkyOONt6MqTSY3d0fE92z6w4t3xGuU3GtOIHGtf88ZKRkRc1SEXhdcO47LqBFmROvPEpn5qUWsf
Kn6AIUcUeXaCaWebU6vMRZbCLATtuG2pvhKwAUjf1CBku0ezSxzCO8rPdI/eQPTuiPI05lg4wXos
OfnhD6TYaDnRBzQ5p2K4tEHx8sFt9wpUEpeuuCeNr2ecED2eyKQfRy0izeoLyDRbwn1jPU6qsdcq
tKY2f/TgwVzY6LlUoC8NjafJjy2nom8h5CWfNPosEEf2ncqRTo0JjGoZEbMbKyXx8492EMmzVXRM
ybLbvab1mqsgE6HaRUL2vgSF+Z4vNHRvyM3zIMKpDQfdjTcV28UZbwYp2yqZYJCVu6z/l+ieBk7+
yLoqPCgSy54pMBbOI0exjEzA1N+G4XIYMtMsKGmqRUAx3HFIwpH+NYv46RNs4JM71WPqEbUkbbmZ
r1mjlHufyQEedC8CinoSaBY+vL+DSW5ZSpa3oQK+cwYFy0dVD/7FkqQ1O+LGYFNE0yeiRCJA249d
GakAVkJSG5ZYtttVTZSkRUwneHmRkPTNwZZlIj/ezjONs4H/1HhL3CEVyY0KXp17zYMAYaSM263Z
fE6rnBLzE/Cb+r8MFmCfw0gHO+2TgjDs61ygS2+1UaqSlhgy+DCmiSNAPvi0wJmDg2z8lCJO6UgR
0PTqUlxa/rUQQEUYdGy19INKKaQxJoe1cIKXu7c2G1V0VzFU+5oIKsU/IASExUIXCtcQ4GiqQfcS
n3UhY6IMzGleDiaDzYjYFuCMyD7z/GIsRDyYis0y+yhJNSWpEBKLqXSdvirYSdhOORHgQmdvQIix
FRGCkbNIGj1sFh9u4J+iLqud7t+bngvUjP9kE0ANIVkcKcmYQNvY1TWofoFnkt59SFXUne+wkUIU
xUy3ufnNl9IDbd5P4/Z6Vm4C6m3NQPBsV4PzoNWmX7PsJySnfAYFCu5Xqei541PImOZ0e7TsLAuV
l34ZRxcbA2QmJniWwCEJuKtb1gHG5k8z/T6+ESKag4/5+DqQJd+2Yyr+J3b376n7QID+jrE8DpCx
Gr9LCRzZfGvgwuZZZLLQysw306+OZD0kfyT18EJBDH9IT6BCcfYBg4GWK5usJlzG7jZMm7VcQesa
MqqVxFVMC/wSR9IxfBHVDALguc01RJ/6lRveJqxeRw/RQy3RRtOPWLOYzqIxBmzvY2mTdVJE3J1E
IFOwXOEwOMUUqEGXUZPV+hyfVImeLNVFqqFy5etkTtuiGl+q7aG3a/1i7YvXsWp2tZYUbWzRiN5O
JkJbGCj0xhckXAu/Y3If0MGhypWlKzDJjnlJaVlMquHOpglgHpO24jGpZuxTwQOx5RzPk7beGqIh
rlmJB7nvK4oZSqBXs16HnBeUXW4nh/Wv9BUgAv/nnsHeqvIg/462aocdQCl+LDK7TwyUsN78SzEY
dCrPSaIqyCxeDCznnDujc58WxOUUSnLhESd8+OaVZeCcuDScmcUy3x9bZR7gWjNSmSyZjkKWln4I
xP/8dXyctVopPnd2qG/Apa7Y5IVx6qoNS9JsJOrduULAnFKkIeoLeBtmYHiVgBnB4yhDgbjj/mU4
gcY8KeuWCBIzowbYpJFnUYtLu13LXz6qNqUyyOumF9UKF6ArbkSRjHGd/ZSvGFyblbdMSVDpND+D
Xe5z1/iKGmUGcr4W2AT+obDZj6BLo7E7yFk3x05kJP9Mm/RyfRn/VIAzLs8+b4nLyDikz9h7+Zky
T4ua3+aVJ6ivQZ1+182D2h9YNxqUAZSCCxH5Rm6w8wVacGGOgZfMpSd79S6SHUbFN6kuZrsd3CJ/
SGFz64kPC9FQl+XzKlTxudRtKZRCMb/KPZo7+e8LvNAR9ZOzcIpof6iUBHp3s0+t6pwVfO+3GO+2
QSFBHa+s1vGlM63qv0OfSJLSVabRE0fz8WvaPYvfS0xKPVyjTfgSSVOBcr5C70VoLRAjn/cauDb6
o7P1/8r9pdkwmCh7RQHgisKkMMACXAbgWTGrST213+XIDDLRux39GtCkrElnmHkimB2NQainMCOM
Ns6BRlhYOr+LcM8tP5J+3ulY89i2sheKS8KKGQWYEu4/aZb/DcESIQqmh8L/6x8TT4YCDRHkYRXd
ZfZxpW72TSXds8u04uaYwIe1iPpzZlGL8RkX+G/daZ3QgoUnoAZAivnazZNQsbCO8DVEuywmRonM
MhjSix/j6xbHat65ywY9BpsfyVQi0dm9HIXd20p7B8kJ8bnAm3clccL9jOFrxmoeHOO2kAWkZH9w
0nEeMxfWVIfwXNSRBs9J0IJyYow+JoNpCfUtXh3Uf/MIfnfxl6pPCQ7W60IKEpshY2yQWpZZB0Af
q1R6Dnnv2esQJc7ccXeJc1Z2CQVWNSbJpmXP4jhBOBoLziJuu/y1MSVN5Mtbw4ShyOdUNkFLqXLn
jegdYF7m6p8FcVT9USgqBT3INujbNSGBDaIvSD7mKGHOEAe1pKulODXjOTz/NfiP8dBQynWLSbwf
ZJ7ymo2ztyFq4as7MkW4vv93DQmBXgAeVqv9ZS85xLSxV25taMqEjNTwZ15HCBlWDBGskkBO/jud
verDa0ScqkmmE75IMzN0LFvw7U1OqhwK6Pyz8y84pM95F6xRIhmKtvPzlUNEMO6jsM+AFi3eS6WH
kLpXUuNPAqpw06JoxV0h+fLCwHl6CQu0Dfb+gtYzLjcwlLWpuSJLROhKIkKmeYegig6T/TDjxKwQ
SWTn1xXMJJ206gk62DzMqteuGgXTVm+qPdn/+YNCWl9JqTrm51b7zPD/SW18HnHvzHtHnI0eYvBc
uTWCMqmHRIA7KtCl37k53fDKQY4rzGyFf8BDJklZ+Y7JMhXko3P9MkUsHDgH3FQ9mJQaHKq00tN7
r5Q/cJNa3H/fhV1qgyJS8Ix43LU6hvcPrBOroT9PxyQWRoJ+Fyfe+ZsqX4avzDofdERgTV+kqmuA
04XKZh49E03OWSXiQ/RGZcBr0w3L/lUMpi+ofFT9YfewF4YuOwOV9MorREbqv4z0UOUgnPhnWJ8L
8/3RQKzSMzJO93znrBR0NaLRIE5n3thv5B2gtQdhoYTQy8qatvQwl3pXPpwrJDavxvV4qbSegYIg
Tmz/fr3cxhTfQRRaCgcT1a66CWMnqzBNvYnC5HBit4GISxyhS34/sLiTPoyopt43fBEy8++I8l/T
18jJBjXWhqZj9za0XG9UsaL84eZ8bAdqAe36wpJLPL7hDWsQujUw7mlHGvhBPJVapuIqj3G7JoFr
N7k2Zupf1huw3YXCJLlaGl8m9RfhqIsnFTDA/0jS5UYkju/dJDnwoHtNLunWP0B2PzjS7xGMUKjJ
fo5LFrit7AmAWDR2pSpTk3s4th+VNZqDgHDHEFMPdHoCPsongzlYIgxR410N+ts8ci7po6qZfLB6
aHLkDDVM+IljhN7drHTbjC2Ylefgr4BsEUEVhzwCrUQirZyCRib6sWaZivCfO35ksUQRwWuqtmn1
dnyN92dwqdQfBOFz3TwwCB8j5w37dZxfJSsua9rgKECQmw3Jb+v7yc4G5wEIcFzeu2MYJL6N9fEZ
LmGG3XLUylYZBQzlDDs9CfWOdb82AnQjlP3GFVGPX8mXAxkRnVZERZP9QPCYTbLiNJsnj/6dWMK9
/H38ku6rXHu8P3rCo/3kCLi2dKC1yvYkJH008YXEgFiC+EHxAj+4l//HmPGLysLxatCm1iuVINcP
1BVcYqDefHrFHkAe1oU6bNn+H9I+3Kp5VD5MIQS5tUldRnNPWhhvPT9fMQVoy0VmZvluZGQjpwbY
XopzJSy3uvMtZ3FDPPeT14mM3LcL2Pzik8Hv/12WqEhAzozfJxTEqgTXXBz9D/0U0beqrca2ycFT
irFKeISL0WEnmhZDd+nJ38hhtAE49Ap0sGrrUhCd/2Fsw9/nj5q35OoIKbshdiHMSJ/+KkqelEuA
SMY/pw6EbLsJmieSWbUfWa1d7aoRWPlDvP7aL5CcgRxObggKJZlmWYWTcbFsDsqk2OWPGgPti4IB
sveptOzgJ2qnEFLG7iBQf5Zz8fu+2VEwlmkkNC/7xhVrHQdE8Naozo+4V0adMcYbHq8ZDjt9Alkh
QTO0qPX5jp1TXS0Vg+5mgbu4P9aUYhPWnzx9mBpErjFlIWu6GQB8QC8dWQrzVwlSwWZda7XJPmel
nttA0CcDsJv2KvWE3zzTR9dH3TpQozVGBLKS9YZJUJOz9lJ9c9tcFNmpDMS/k9g1uAKQt3o0dxns
FA7VA0JJLRlCparSmYh0WDVe07g7LUqGWcGSaOXg+Ou945T3wnGpx7yUpd7Ctaqw2fMfL2wgwVKl
7WRiwg7YZ8pi5ab02mXI7cof2b+GiYDJR68e9v+o0ODbVRiMpSDP8qiTEXPdsymWN4ObV0kodW2M
eHZ/OJ0sOZnIElJ9X4tkwy4QGOHmw5Alcg5dlW0KAG8WW3qVnuWaB53yaxHXovIi7nQDZ0cQuxQS
LKOBz7sWvlT7hckwjUPhK1kGZki9Y0S8I0LPxnvLS+2W4o/ANZZ/wYoeb5grPYXb2RR49mXwc8Z7
WhabBeuSAwlx9H1xLwsaXKzy1ioMoxYi9xjYxB9BS0NY8xjFHLGtCDxjhARsiY9F4d9Yh0N4c0YD
AvcvxuOUrZTAl2SCSz3XWNNteIXJHGKpAHSfebsto6VjsNmnU4blsXQoZVgESvRYbk5afKnypkY5
bmkOK0bTpx5mwbo4Jg4re/FDhvG2F+8sxGUwEiL8EuK26NzxFUbZh/DF6o7uCinSSjuFA7uZLDJQ
Wy+YNBvFUZu/l/dY8Z5AAjoEoDeZtUXUUjaoOlM5OCRrg0nyzQJmTw4+k7lMQnNITom8/1pfOuto
z43WlPTXxlLwP9Yujqje3WliruyUtEo+aXHyzOfWqa9BsuyXP+tvWNIa5u8ts5+1e/Pcv7lXHh5v
3VGXpdC0eP+MiHq5RJy/g7zzUpCUw2vgnPIb4OyqDRjS32A+Rzi8fMnmdscoSm2MDYnBRci2wmaR
fw7SAL0sBbVGrbXS23iAx/SYShrWJLIu7G9M3oOOwLFxmjCIM9mqFXeL1lbuV84JIssLAiEJuAiP
suvvCGufAdnINheAdhMaKngbdCpWGm7+OGabA15CS6zMjXU1b6zrprR3rXps481JSxvMoQzYp3sS
yWIYlMesmoBd5fwGqVjyczNJxYQ7NGkHwtbQbRaYyiqnEWC38fMbC2zBNqAWAX4cDjRBJWUCFdQ/
9Jhr9EVz9NFjvWHbgOQrpt0okDmyEue0spTcxefKNKMEIV+k2WHIukonQG1TOMDdxI8IIyBZlhGK
0ziQTgCRRwWYwssTYQmd4Rs765grKTt9UtWTerONK6q3/n77k7xcaVI93ZwIi2S85pePzEQHevO/
UKfhYpVBLXnCeRYwabzkkM/ekq80A+DAumSUDZM2kqbOVgbMxVHkm7NiP6SytlkfxGiyNsBiL8Mm
jkyH+MgP0ynmA5ad9G962f7mkTH1VwsMbPL/CPrJC3gSNKiTBqpNuVkxv+6IA01xGJalAe5lJIlD
qjpGk4vCDk0EXi8zGHJ9Z/0tKLrHgcGIdZS4pSwfGJr91QceNMuRud/f9cHYRQYhr6xQsF6/DLrn
vO0DVL4kAMAO6wp+ViqkGwJj4n158r0vAixqfTV5wqZ4rTVD+5S9Fr5UvflZF5Shs0Y/XDjgA8UL
3kuoi2sJxZdUvoWOqBiVUknewOsSBMepTr4f+KI8HDFAdZplt+s/revCoc7BaL3R4OT0Zg2+71hw
fBpLws5fkG8QIywZKB1yxWLFFdg6uFPXO+6xFyJwmc6FFfG2z1WMNOGOkzl+Xyq6gyWFmP0MQ3+n
g1peoEM8dklbR5X5/ISU4h/Raz5GYBKn6nMr+FmKxdiCVc1529m/oQDgXqT81NU/2wDsnCp1YH0U
NhBu57d5vKCnOAq42JWsT9qRwSOxC++njJZIVMjx90ceXI2Fb8KIq9aAhQyBNH6A+CcreIYfrQrU
nD8H7kHiWrwtd84xGIwDoeeQFpi6hmx8ekYZdwDhd4cIvtXIEKyu9Vf9Wc6TVDFBVDLoAfJGfZ5m
52bT/qrOPdGN6NjERKh9lEcfJyuziriD1l25GCXbj8Delyf192IJIbUmhqcAGk3Y55xTEQx8kTn8
OZW9rdxCZdxYmHDPrZPlEXiXao/Jiy7XivpQ/2oxzvxkRKtATXWs/tBIWeoe/x50ijw5Y0tUqVMc
qjiy8sPBMqqcW//6toJLHF16KrIVHsn1jjxM8kxFpmNzF/tlbAaXUgHsAwkW/Hm2CvvFJH5TnKfk
G1DIh3/DDXNJeAn0ZIM3RTOmf1Y1jIE8ocm3n5fpmum6dTL7mSt1X7tP8LXCbDd8HI0Tvv4DDLWQ
fyF2IpvEGNFRpZ++Trw/1/jbu4M7c6zltJMmpbwWMJuSQdz2krYJ9K19LzAnu5JzzgMAZFwaBq5q
MERjHUROfHgT++9uA2cc/TrRmSiUyKdelqf3D52S6fMZPdzFhb4iRiPFIAgTizsPfWhYE0wYS3wB
lNM5WCqYmYp42yI8+fvPBoM0JyLDcM8LIpRq3CNg5cDoUnwuzVkMkgwRXJS64NXvoINMFKszPbj2
ZUXMWVygvMXYaiMhj0rNw55MAkWt4q2+Q9/n2HHV05LofT6/ysEc7R3/Owlp1H48QBw8tboG7TVG
Z+RuIILTcJRSYFnwDIHoB9f2gNroGcfo8xiLN9laV05pP6nVjpPXjxIcGUJH+IGUi5K4VPqSuaEv
TMcQm4M3qdZ7/+guiI1ug2duU8hSbeh5+Q10D5qXU5f4ciGUnFwhsYYnNKMS1ctu//w3JhnUFMwp
yBxxJwfNrggtFWQWm+2Za3rGzlF9N95SHuBQkSwsHwFxjemAC/ofCtpa3i4u8GxVyGx/pD+FpFKG
ok+8LS9O+lylt9TSBVEdp/TPK2SCPFSnyLYNhm4Noq6+VwzH1Ru4OvlEIZ9AUyLrkkGc7rYUhaSt
smBY6fYIg4ON80W+u3ecOTjrsr8CMccfUdhBzrGkcFEhJhQx0rRiDHhZyoWXL03ZBSSViXpo932m
BscgQNTmTcrkEaN/ypqXqGcIxGW4pDg1mrH08QnI0NSbj+qg+9vFDGE99CKpKmFelxmCcV7M6YyJ
a20Yc8Ilts7hs7lSXf1WpMUIhu9y9uUjEx57keArgGo35PJS+/YaCOvEWfFHwiYt/Qz2m9ntl33A
cTCquDI9lmFIP0qdA1xnn2en4sbLNadZQop1wghnb8Zq5n7sT++kkH2TJvU46KE0tYEni+erKHxw
aI96aqqAgcNNjjYDechIRFase85LrW5UDw2evs9ZauFfREsGh//nUCQJXt6/iivCYn1hhVfiAtvA
hiN9s56jCvJj3qAV9ugKkFcgWDgsql4/Bdhf38Y4N7noQiUHjNtlbO5PeOQDvbhbMq/VavKoqZV5
tV9FBfgkel/KnZWHG7X2bZ9EKZODsH8DbenZ1Xb+acBhbNsOIOTv/Cp1PKIBmZNsZ315Wa/Zgqgk
GOpm13nQQiypuJTLiclYWNXO2hpFDaL4vATO0neHiI42lNJO/vsEDUvRNblKGiYjKJta+sbiNltu
mEfVEb+GBiWSdDbft36zW05wGIE5WF9NG40j8gT5k3yjv/SogQFQYQMvo1/8VZP8FI0Ffhq2wiZs
xekBLyinQxyK0FU2x64zoytb9TYjoTx9v+68CmHr7oQ/hQv+wUxrF/YH5bgKtyVx3oP99arvPzQB
9chC/bBPSabcxHqGEs0DAUI+7HyoI0aNYR6XIrc2L/SX9A/DRTI3JLH/OZnhgu1DeyCwO9rLEqw5
UnITeVGh5zKfD3jy+PEWv8RxpNDR2LTwa6qnd6RyA6UmHyetfN/2DazTasBNFtSXm/4n0lhiscbh
hSYeaG8CwmAwI7m9m2vLW1MiazRCFJ/6Ie+xFsMPUpPLThq+4W9YlFV+nhlDbUSoztY6cmNCd0QW
dpy2y0rdq0OWttG9+GsRiMXIODWNwRhjL0eeSIZyL3GiDs1syaLBasNC6Ddp/ALnzAVmDuddB35D
WT+qLKNCJ7eDkftqxRo6f8EggMcXEMuZ1iUGmzRGTCxOv+c0i+N285Xsd4CFv0PpEmwrw3/w1Eq/
BiyIkk01L20TYjV11VdFU8pjiHtwapCPupR2ZjkZvoKNTp9joGVuartL06GevObhqa4rLQZ70c6B
xLr/q2v9Pl+P0vQAcZYxr/dxzkJoLSpahbzJteNeHh3IGypUdS5gItH9q5+Aqu+Wa8Y2yE4xsNhs
YH6VNPPj+wEhLXUGl8i3ctJBSXJzFx0+4yV0WMLbqQeQmp4UM91LF64Qe9ATsnl6tVEEBVBXSLMf
nVnbEQ6xXUeOClmrOhOKDZ7iZsC9iH/4NYsF5T5wh9PCnDRs3xcoMLjfXfOQRUqvXwtPcHP6Q55M
bXyQ4EbJ9QtO3RVzZmOQczReZ1U8TEnqcCTGnaroxNby5hgYp7SDlutvQgwNnUiooW66LCOmbzKK
uEHAyHyhPbdUyXyDkmPs5zhC0hNlZCW6Mm/CV8qyguf9Orv0VxIxfO3xLjV0pAlZ+NUfxxx5yUVK
a4W7aY/+rmuuPkAl0VWLhJo9P+wletlRCvAvXrmKlDPTp1QVc5kuF4Kmzr5vQYkbvMjE2IJb+EPe
/Upp9WKLLepyf63d9c0lAxWbPBMdgjaCdpZUBh+YucNNgWKFiNadDI5op9aTWu5EQ7ZwynoIMYXf
ygYYBtjjv8yvwIqYfDWsqCVFXdfJ3TzJykd51WdgMqJR7AAikYuZW8ds/JRTPNIeq+7yZV4jf+yX
hgxANYKRCv3WpKLD1rkffzQ//I4APisH17UZYGSC7JyYx5c+h8ofHSL8Vaawf34CWE9Kvb6HLPNY
flN72EZsChWYVUu2BmAC91ja0o5wKytRdbe0ISFq0C0xPDpEo7cA+vH6oRUar/b4lKwDixe31Nrb
XBgKiDFbIX1D3ej6ZudbBt9Dr44sqwIcVXJDFyBNUY4vUl4WaL22KcWL0CP6ZewF7KURmM1RD7kT
zEYMORjO121S8ENH3VUBanwUYs/j6gu+2T2u0OVxRxxmAzeIqs9LgW26YquMUApBhu533Bahu5/a
vzeKvRSk3oUMcLNUNFc9RE38Kk1naXv2b+SAOT50i0azGYJR0x+DMAcC67sxkc/AF3VooMVGW1uT
IhpVORgATDrHkSo8PXTiBBp6WUisLvpyrjfi0uPh1cwp1LgbPy0S3tXIsjan7SHd8rusd0NCTvrU
J08lOfyuQf4VmP63jFzjBjkiOAtWP1mR4qONDZfUyXagprtyzbOf+hKftcrHhBXvgQ3AavRsBA6A
Iun85XtXKdDYNfQbjGAli62l1GK1EkToBdB9P+XZcLb0+VRzc4kMJA/9V7RZewvBViPOi9iK8YkB
nIy/6Y3TwbSzTXvLwD4g6OvZl7hW4wd6N2suu/WT5gVnnKjv3xkpavSfJCdFgX82AiQGgjbKLpx+
RtBElXtqP5YpapWbqDjtNo/iO1z8xJew7n2AyqP4Jo215k8Y7d2K/k84gmi50jOtCzPRQX67A63N
vV/5KwlM+sOwMyemrn677TKO1UXKb3HPPV3KbyaVT6ov7mcrDXC7+ImNXTyteqndznro6Mv3a6eZ
ND/uR7pj2kGRL3N9mszq4dsRKCZTPzf4l1NPIViLZVaFKongtH0d1W4O7J1vBVIDmDakvjcptOvp
8lW3deQ0CGadjoea+xhh/6ksvqLzlWMlgnj1IOq78OVkTdW5SJB4giU874fCmrAgF/8KSq+hIgJw
btZwbNOi1BNi98V6gy3ld/iJZ5Po46pWD2JExGyB8CQxf+ls8wCqC7Xj2YvzYw+a7utauIKZTsat
Eex/XSGKpUpBQ6iTLW66C1H9MACwLCHp6t6845Ip7hm7W1CaXJzXTwx5keAW+4h/2SjwW6bKQUB6
5wEzWAAKK9rnC09nyJHTj5Hbfdq5tUY+33ikDbjKLqs4ejDJhihJft+GxwOW/z+XWCtMdL5ccSj0
21BHFHCCXw+shbVwaj5swBBMjHMMKN+JNuAkg+oWMzPZQwNrmxY/3NOV6HW5Ae0ZRqrHX+Nvkot1
uXiWWWlZWfb3eEsSH2BnbNxUBMiQe/H2XIHpRtqiDH/ttNbDodVCyi/W/hFxMut8gi5FUwV6Nqa3
E1jpsbzYrNczIumuR4TNOo++JfPip4dIoMNtAG4SjOSGlXS1U30Xppgs6Giw7diZRijgv2dZiWvn
ZiY7jIf+/R2p4orLqZszcUbvK31bsQ1DG6uOxCQcDl2WACRU94m2Mls8YeOVJlx7kOuiN2nUumyx
0U7wuLVP3phTy4A15ricWl79IIgwPeyW+eAc87JaVTB/2HlYRiW0ZKo1JmHTmVEUOBKCysuXhqgf
7czKljOunVSmYOcMY6kdW0d76jxmLBz5TqSTRO1F9BPQNrG5iQhsvl3vsuzF5ebe8M4SThsWca/m
qtiEciWaCOXpy73RHIKkyxyapZO3KoOsz+RQ+PmWbeJBbFHW10K8PIyY4yg9Lc+ktS/AbtxfFKC4
jrU1d7npe06Joy32N5zOJQhD4innGzRn4GoXRfVVC83614Eu7icmI+1q2WxUfP5gO/rvYukzs+Dt
X2HI9kvAjYC53LmfOInlNevtfSZpJGkdFtU2uueh9Ki4fOT2trKX4PG9o259040j5ltOXHqWYcs+
29AgJhmTvM7rxxqNUGl64FFPp0N5JXyPhlvryQeDHyM3DZ7UttbsOjiqyNNL1unHP6Gw8T/bWcRx
KaVY18oHojcYbV+Z82GI49GXatiiYhl+PZR41tSu2P51AFUqIqi5RfKDy5/vfGy0Ao2Qi8exl/0q
HAny6YEwq8rSZZAav8XOrqbBB/RxjALyjkoRHsTgjZw+NWpxMFj7Y5We2YDlxY9l73Oc0ZGsL/Gg
0hbUJuhz4MmCXsQl7N38tRBtn2vDzz5/NLefaDRuA+Ysvba3M79BhEjkcWtzwHw7TBVumaWDTgf4
Q2CaqBcbqij4QiQHz/ZD+Ia2PAdrFIYWd+ac1F686yQPHPTbI1EI4N6Xe7z/7Lu0L19W6WHuhwpC
l/kNf5FJHvUlx4b6l9lokfk4TOzE9Q5Cjiv4F1gIEh5+WXxGV3OXGLQNYII6Bf+lsNtu2RLSKzq1
PW1lZ4KY4//TMNDAYP9MaBpgOYTr67Y96uVxPIT11wO3Rg0IN5MHWVgzW+XvavZWF/c0RdZkJgxX
IHphP8X+Lvc7AaQSBVsW8rk7GBuGi4p5Tb5c3kDxAKwmNprA6fSBhoo9oEY6CnVW5e4i66QpkP8v
nfW1sFVGK3nKx1cMMw8oBuqSqELq4l+BGr8VRO30BgmU7c0F7DWRRDpPgDhdvh7HQuBgXhoqnglY
ofSwv3h1oXg/tdKc67+pWOPBWr3DiiuOXZTRQAWggHrFSJfM7LT5ySfAJv0VbRt8Oc/FeQR/0+5n
vOKudV+q18iB7+vAVZPNVgLIy+Etok0JTW2X9rOd10pLlnWv8wDV9V9+uYY2kJhPL+3Ze+1OGvG0
cZA8pLgRqn2GV/aregzQ8sn0oFNQtRj5r2CLNiufDtSrOtA5QUeco/M/svBsLhYP6vfQ+aphbDLF
VSJNOuBPzSXgKOtz2i95L7dHljtCCR52O0x6iCH0WvVNuIGTohTNDi4nmaffXoZ07s/YM48algTn
hYsJ56jGEODKXZIspA2FOUW/WqedvUn3rKjBoHauIzSbqHX7M3kWgHVic6O94fo2u39YPtuBVRlQ
TFhJklEbkuKQxC/x6l+lUQpuaZfpgmK4LcpPLiNkuYD2C3uIowdHI3XdlM3G9k9EOuiTo8nluR1x
hdKsqPR/a9BsOrz9YvpJFIJGcGnt7zIa/an4R+h+B9csvfO+xC2EjWPEuwOjPVmVCyY8DGqgkHIL
UN6HFhQnU0OOXXa4RRCK8dbmkIP6HY270rb8JckfB4ualUKytQt8Z1wxCln8k7jrapNIH89IGc1x
sC2814eeo5KmuO3TOF0SB29rElvkRjYJmSNUEVaNezetRBL+ZgKGyqWF8ojgeXstZs27lHSfHlqe
v/AxtwLPMXsao5Co22kLd/ZqDUz9f8eA/GVRv1P4jVnYzS+y5A2bJsO86N4ROd90uE0W4pzwppgq
g7AUVIVR1wKNa0Vt96j4Bpb+G7O3+hrpUxduwj1C3g0q2ZsOGsP/oF3fZfvLjM0GHjbvBQSR9RxR
lXAQqJReAUWg3CVnRVld6GSmDkqPSmvmNNLr2hLIus4UCXZQ4i8b6j+Nv+sGZAwbb3tkkmmH7JB4
mm5z1HTSUbxiCceXqjOhxpFg/o8T5/ROtIo9FSJS5wA78n7GTRZ8AGbuS0nzjF4xi86kYrSo35xK
K73uXK6+rIRLf7DmSwdQ/v07F8GfFYcfCRBmu2EODpXfKXdu1ZQjaY3OBuJTQVYGV/2XUKg8fFr6
fzDyB8eGwHoS+TMjfh23eYBCo8G+nslggAQ8koP5qyQeeM4twVqCRQpFKTO03DsMkd/D6JJDI4by
xqO27y5uPEjbNPWUEKozl8tVemw38TKcTBVX56uj8rJqYaLBKVYirngqFXRnKSv2wVdhG1zPNl/T
OgcZCaHYfyq8DlJzSRPXX7euLFpYyO/PeRAKNGIVkgSZwkqVX+a/FKqditHQBFjWKFaoheiSlWyN
WRdqMP2DHcyUUXFZhHAIu24kVpB6mqPkZglqR4+rgu6ExJkaTVO+bz91uI3E52YLNZd7K3x3m5MA
xEbMN9PapJn2RIuuyumlFdsHZgvs8QuknZpwWxwPa+vjw5AzRaw2xuVIm6QbOV7Inb0GwD4Qzm0k
j5Xc94NjKB9ZqBBXpX8IGEi9iyKIl8CR1Kw5StUQs9skdLq5PDVK+hURlpYZFAlg5p2Z0wlVuWTF
3X7e/kjRWG3NJAUU4wX031UL64zYID1r8NJsI5p8ALpRpxDrjViH8cEFctLZqurZWNrmlJGEafgl
NdHlvmGmUJhOR/ObFQ9Vm2VaAWlRNeBTickQBGTqvvEPowvzQjWoAqSjeD3hfuBGccCOT+WvbzYw
9ialIDkU5Cb0/piQC2psrgoR9TMQ/yJP/K4TRjoB6nfdz3vwLP1dN2VLG1FKbbqmBePgJvdpn96K
mbB4mT3YPtDcBxcYewQ7qF1o08sEwR0ByZYR09sIh4eWKX0JMxYxEGL+AJ9SovSxY69gjxweBCNB
q+eUqeW9s91VGlQziqDLh9Vpgp644GOpaAAxG/dJKQnDQlYYSu0aAyOtygtC/ZXUuAtk+cah2Pr3
syv41XBz2hi7TF3RSX8iVrZzrUZ48urWscMM95wZ7yjVxYU62eUpS/VooxMIpgD+Jslhn4KHx7nd
iYKkRCw6xFMg4TEYQYPVgLYc3LeO+Jj8XGefKp1oVT11yQvwXC9EGylNm7Jn5LjZEUHCDzRDJy2r
7qT/BevJXN8NAymMec4tpJfWrT/5FS1r+0AxRwov6CLulxJZ1jIQNjVmmD1WMhy737yilT9PMsI3
soDy8GTUQ11GFqHAJnBwD7eRanatQYMiYNy8Xz2j41C0/nGl1zq6TYlSD+ewdS9UeyTHqXxeHBOh
jTlnwRJfT2CXTojh/U+hjpGlfiRp+OsOzxA2Ihiu8vvBYrN/mfD+5FGO3pvPHD144ZK1LXSObCS4
dcSRt1uWYyGb+2Y9agLAwv0vsxNgzlH6ieeVky70hTPuf/w0nwmHHX8PfdWJajs01dp5xlozkt0m
xczhdEJ/GTdJI4rQRtCfXJcuT7vQobph5gB8PQrh3nsS/A8XWkATM15+nzAsGpnWwKuTHqW0PfOG
Vck946PPHbofoK77kLLe1whSgJRgB+MzFnJh/lWV9+TSuqWJNYdUd3/1ZqJFfJp7Aw/+3QMduuMd
du74m5mmeseWVMRTA1AxBLeGZtTuPMU22ATW3sceYTWRLmoATLrGp4Y3n0E0JWKqSnOD1wisaMUR
MG8HJGnYpRQXf7Efraq5Evt5sfBh+RA3XEzY9bdLYE1TISoD42yNOx+Tghx8IOJLnUXnvT+G1A0j
RB8tmVQ2jX6a/f41umx8SpjPzscV1uZoMU5nx3cAkd/f3zFNnwAMlMsvcbmvb/SmjdAGPtWGmlae
SpQuXKmQSJvOUSOuOfqJ7fWP+Jc+Pj/4lKeC72fPw+5ZP/sweaHhV+qX3rVaperfJXzzPWM5P6G/
Z6c9q4Vp6VUJKPwF+gnLcEuzaHA9yC8D3c6bnjZAcMUHHqbJxTyRERKpqBbSdvZauUpnNLDkfMKA
sgNwNjKDF5rOp7O7pax/yrJbZmSHVgfxZETcaGsS57a+A7AZ9RCg11Ax+5lNkk2VQDxaVJS6x/oL
OLmqmPFBgZy0x00WkF5l/VaHQxwK6KxSCYe3AWuPANQpcYWR+NuEAiM3D805U8rBLtlDxXyNGfgo
f3Y7vZ3SefRVDAUTVOGpmdyPmhlLflIwIfKlyCBXcOuS6K+0O51QF55Gn9nE9WODWB2bE20tm/f4
zcBqi4fTss8ittjDlYLbAFgezFf91n93HrlXDHk5W8iEymDto9JMxErXEg1HfiQtpGkY090rJvxz
goq+zWNeIM28TI0p3sYMNSotxcBlNgY4J8rn264JMAXRZXaTZNcYssszd3W/3V/+jd7TaC30IxEb
rjRK1Elf45q1MsTHpGRjTLOTdMNtU50hgSeJK92Y8g625HS3MrxIeX3LGKD0T8Ime2f98MHPu5cx
m+yKAqoi0dWP3PgJA4gmC07VIbG39U9uYuHBp9YwKvs42RpHeGGv3oXw9nClse4z3SqsAAc+tVaP
1b1/oFZaAuySnsmpU3X5iGiFdJCenAoemFxmSmutKcBcuaftrdRtGCCYeQ44CuFcBszE/Sv8pJjz
CCnftIF9EKPftxf2STm8OkdaasgnRv6a5TmeXC0swEgqoqoF0MXhROJcEYkMOpXfV4Z0Ayx4JSod
Rxt7IaT56O2vkZ73JlP1m8bHUOVz1c5Ai/7NTHlWbd0AhjZzIXvvy1w3sACLJigRH/7lEXgMW5pR
/1IY+8kmOIfoy5UfxvxM7GSihfxoHAM8EK1RUM/0RG/5pN/rqLdkyU4lVFMZBpx86U1jfmmdsEvZ
aLmaZQIuiQUDa/zd7YoMLkf0321iuUH/aDzpoqKqOgGwag8K8kpK7nvYq26EulubO8qlGiz/c9fK
6yRMCfGlsZuPMOJKVYdeRwy4UFA9FWEWd4E7lgnCHQK0MKHv2I0oDlNAJqlrPEY8aEiwLrbOY4LY
Hvjv6yDuv3UNmhKwtgr4r8EKIYyqYZwkH02kRxg1gNwG5X+zyAZwZH3cc5NiHSsDX1gjBQqwew2M
6I49gOXTkJfX5JGihhDWm7uB6iKkrveX8/TNUygKNgboTM8Jtz8wshPRwtCgaOJN0JOBuM96Yida
64SrtdnhimKr9EgX547oh5MTaZpBVvrTyExlBq+A71rzX/J+NhHReLTFPH8mnW8ftU4UakXPyNWU
LG8J40AiZ2K2vahRA4gwHhzNOh71+OjfMfIqz2dqrS1scx4OIDTiBDJaMYiYvyHDA5yekXuSqjCm
HZv+J3t767z/JX7HW5s4ijevmbfjWEIBSnLwCxRGRPRr8mlUDYrXK1sLtLEZkxu8oT79gcynC1ls
c0T4eo0NITq4DcmUXKiACKVId67JXQnbhfrFCajaICmVwGyFnxuJEabpvcn5e1Nza3rFt66vpXVz
bX/lZbO2eAFhtxdgp/6WZEXpNlqk7W8bzNfsaZs+5s5rrLp9N3nNIxtrfGcUQQmwMdm/4lbcXIh8
L8cR0hbs2oOd4hJ2T1BsKSVaEYyzG1+h+0HIuNaxbiidSy975n5OmbG2x1AOUiyIMPcdjtq+MO0t
j9u15mf7t8hUggNIbriKd1BwNsFzaEqjCVLUEwqbU5A7Y8OL/agVrYjCMG/MYLv14Uug9GjTa388
SzgrqFgJXHemwrO+r8Zd+qRvJRqxHPg4VZBwc6m5l7PsbEOAatBGIsL39wPaww/GnQkcApaL45xo
kX3sjJHZOwBRbd+SLQqOkJeXSAdnfvj6X93iow7uiadtRqa1seAZMXAbJmdujsNwgCuivSjEWC0m
IEdQIXGquztVN9LYtrA9RgYpn2DS2+eoEd4urT46OdWElIzV7xeELWDuI8sJ1319ykjVkhrFxpbU
b6TrQPKLAYSPf9vrWtdb9sLYSfn4lrQ9Fblg2oAi26l2TnEb1y7WTbvoD0ZOzCTEqw/wpJ6GCj/x
w7jT4mTww6P0Wg2OuwtOmdFwD7BsEu09ZN0huB3K10lgrIcybfuUL7ESfX6DTC78MMQvqOaVL5b+
rCozul/g+JfgKjoK2SJBxtlNXaDO2NJOyFRnCJijMNLsARHwUTTo9FGA7a02SUkxC4wPyziZrBUL
Sp24PXKRfeqWb2YihRMzSLzVtkUJu1n48b4OD1H5LxxI0ffZjYK/oZO3/qzAl8fHyDZio7ldFCzR
W4kl3EPlSMwfdcgUlorF10LSXd/m3IBU/PC0E3CHtOztYMa1ucAF4MFJXtS6obq32Oksi8IeNbW1
zzbLlPhHFAp0Mm3+WKthsNuElNFIIxyYZ9bgj62KHDJMXuUvVkOJ4ggQlbYwQqFak3/GyePmJZ4D
KAaB6LTRIxmHK7UFFEETEXBUestMldICkvelDSqZlZT5fBiLUbQFZoJ1GiJNtKfm3ja86AbQgVsz
BQ3iutiLgg/t3t8Fo9FRe5qUl3e5VHFF08Cqi4O8R9BNdhD5/Rb/gAo8J/qzu1kRkSWvHHqUVaRI
8zNmk6YGxV6h0PMnVuHQDv5K+OdVPN3cCc/9na9OwP1efACNxY4xfjH565DjL/vngo1jG8P4vvMF
9ZvqdBcuL5m/713TshxqzAYOpYpz5v7ZMyX73Jls6SdeOgHOdFrUZSwbUCCKyFi1baabLzlKwdud
2O6DdI+ihiy3oY51+Ck7ZYqNMHuZy1MZ50YdS2v6SnsEXIWniroP6VG89V2bbruhNsqk/kGAEXN4
rxuON8Szv+8aDFdPPljKCq04iilgVP/Xlx7hMuJfbzjflqGauy40Etjc4bt4klCTnXNEf8+p8yJB
gGz5OZ3LbqirpVi8TWTH0sHhNmgcyxQ6ZGNOcXmYaaiPi/ghlq5Eco1wriGfIJnNQJs8A95WALUt
JDlKLSGyRLV7Q533RcK9TWIfYH7kSgR0Hh/iQ4f1bFQOnK54fFfAICxLiudVKr6199pNH5TKWaQZ
ZftjkW+5z2onB1ZyZMC22/8BObHpLK3H1GpMFgBQwiZZ9SXPiyqh2JiDZJUH8B49ErMJQdJ4io8l
/IGfu6m8ukpFTSOu3DDyb4BeHA9PwE8Mpbt+qPk5O7xdVmJpWtc+y2rdQjRL7WmanqNeMNhnwQmJ
FWQfKUvWrZX54IXP1jUwwdwYZ1G7Vy+TZLT7lmDrd1sAyIM0kwQo/5vPo9Io56epDMSUbq+tl0AE
3p/Aw49veBm1QN8bjBiJPVoIVFDvHkBaoU/c4Z3mqVSjnNkEYJW6fKdgTIVZ+SkkxA3rL4g1DxYA
IExBQdVm7l20Ej7+m4GQHeDSyxAFbIDXQiR5m+EqhG2Zdz8op2lH8ufcohxYAS3+5LSNsRVeHmuP
6aG5l7KhnZ3k3Kui1O8aO8JmS/EprZkoSrtL0iEZFap83pbFGCch97Zr1ePPkC2JKbooDNyEO2Jd
hmczTU0K3WlCcqOYebNp9ejSqWlgNMSJu2RrCCKeLdeFC2xf1XGDJ84VrMDzQEfEZhypZwhDJLQu
Fpl6WwU3FkIjfR8Gy90w0TkVnG2JEDSyTHnP8cQlJ9CUeOjt1FO2HVpJHOLlHNSNaxsDbtUuTh5S
o8e3Pkh1mxsqFHOxwsxyl9syLdC1LS2NqxnvoxH/zpeHKDwjBFPmk9fzAnEOpIo/8lV/jauLKyyy
Fdc2mMivM543+9+1WXuxVkOxPVT9vhlQwnoISo2E8ykDjt3RLhVIm0nvd70v/hJMOdqroQaNW1GU
0bBK3rD+9ziUFVbYPASlYtUGIdGntyqxBATHZzlaOO1wmaYRd+i2YWlvJ8wEW3dHoG5AjbmnI7QC
zkX/C0HinFsbTQokRCGXAKHjxqsFFfw5qtFIddtzQBH1K78j5Jx0Vp2EJQgabE4oM//VfMaHgKAs
0n7IFRyUP797PZa50FsdnKh9Pmn1db1x5Fr5o7fA8IBTDT2huH3mbeTm1YHodpy/H/AaCdn8l9en
EJ8hlQhy+cfq1Q1ob3vAEF/6mmjj+PLXr5lMrnVRLrdNu9DnvffGQdxYNuZLjMnidHWBqrr8t0MF
jC2/mTmb9PM+6Bj9q7QWHNuTdnKQE3KgvxUGrSfbM/bVbeH3mx8roC7GjfdDIKAmIFZDbAPQKu9c
aL7aTxEWNTa/B6GZ+PpDzyGN+23A2B+HUbZQ2p8oyKCNBQ+MtN1SXZSC/SQ9NsbsRBe+cS7+zQ/O
RgiXfpb2kZgBg/TsBxcfopKZO3gvN1F/y5XwerD4c9ncuos7oc0arxGcx0igfTN2qHIQZvCJCXrE
w8JJI9OAHDOe745+TbsdoCu3mWNHff5fwHNQQ2Gvo/BnPKtUD7IzoECiEcGitH+fFUodHR5CSdyl
hEaS/TSKGLyWsyVUjz4mun9NyjdYZ68pkNxfs5YgkbB0ityww3Q9aBXzLaO3NcH+FKYZEhkHh3F2
miiiRSOnm1CvXS8PcCYLt6xweTIIwVwgcjXHK40Bh+I/BSv83BAspOfFMCT/0p3Du5Fj+BybTbaF
aavP4KxFjwxlLpzk81gmwt+f8zBAdAAC0jaX6BkaeAmzuJkpTCksjNLeiwdbM773xIvSwx5IWw0u
+DUNsXomFCoYTwbCqe1ce6K8PF4lwBAPCCxfUcHatGFy9XLXDipn9h7Phw+nlhl5h2zC+GSffGbx
DgpFBU0ZnoXP308ROrxdDMwPdjJYIG69jntqQZhLLkzS3DPQnqJ1S49LuVPmkbMnfghsmokRNkVH
FB2FHouU3qAsMVDwn2Z0XG2Pb/o4azPYD7IgPrYICm+5iT/zyrUuunkS2EdAydf0T7juIpuSiAmg
jMEHOcsY4E7lGbpK33MHNyeKmdBi/1E0dr6E8PiRblkvppWfo54BFYQbh/ipqCegllnIVsKdmqE7
2EdxHj/DPq3rqKzbLtggptQH7P3go7y2G16HJNDCp2ljCl9SBJkWZhdeW8FfCBL5pquqCbkXyTS8
XRYTFk6jqilPHLEy4y6BeF4FGU7I+nzpqzgugkJqNnKKTzosQjf7keqMerKRTIdOwVic8bRzx5yi
4t+hgN1/ObBKipFRX1B8ZgIDFnUUYHlGf840MzUcTD8UmhO8OAnjTopkYtv0qJjaulEziQi1Ua01
m5WtgHFcKO/6TuaxiyxScewBb3ybDSj7jpvrI1eeDEQy54ibyN/ynBEJDckNp4YeHA5dLZYzSkKH
LBd0rzoInEyjAXtglKidFf/J9b5DYmWHwo+xRYePu6ey65SykJX6hCJwhJwBn5V1IoRtMy+rRmHk
cUK6SiENx71/b285KZcPx20PQPlBmDf4KOfkiYwRJoaOKlln/KRb/bnFhNLpPmT5VjIzfFXIt2ED
Utoxhc6TTmMQYH5m94ihCTYT9lYuU1dA6EIj4YtHdHGRtkINx3jiSCAUK3aMECE2p+R8XjMl58Vh
+zbo5nMvbnG480TZaMytwb8cU9RoTwEWUYDEVdmauIIZRhJaQqUNg5swfb7wQ2Gz9FblM4jb3uPg
DYdaQPMjhwIv9m3QY90Bjb/PszdaD8MiFeLbncI2at159zzh3b8Owih432x7tF9gccwzEYSV+XNS
wAmdGA974TYw6PUuaUufvrCS8RmjQ4O7RITriun3PkP/eMnhnHomi9esDPzefFl+uP7cSdWaazkF
5ZQA6tDEuj72H2ryGTRbrj4uWIsE+khxhgq1IDken0HM5Z7X3Kznn/V/D2k2pD/RyGIljlV5T8n3
22u8yIMze7/Ko9h4O4OVZoo4XVfLXBysNo13pTWfftw3I3k0LwiwZqixzqqOduAkTSPHZ0UTB35h
/6wRv0jdvQHDGz2yKcghIjIswqHiGVqhP5HODFvm9b+HynKS1KNLPyfwjdzcLU/Mf/lI4dnJJALu
84+TyRtGgPOKEA+zvUrwWox8Po7S3m5HzGQDHpuIk1GPmNnrQgE+aybVHE4ABIBffdYvSntvfsID
fGmZU58fAJIbBXOTya30tqtbZ96va0cID3FnC0rZ01B+QJPbL4asw2Dc62dN3WG2N/SwExvNVwsf
cz4tJf9auBG7XO69FIuGQS2oZ2SmXTZr0TyJ9Lss5yo49Xn8m8pzeVasdmX/xdPeTXYZvnobVg3j
KO4HfPKkMW722Y2lOGZxkKPBkcdtGk6Sdb7rapVfHrenz2X7X8fVO4Gr97ZBhP7ojB3NUyfKwzZF
/1eZR5ciEpoL+KfaVkhHzTPa5yp/gLtq1TSnHOyPK5EbAyvAGpwTtSkRv2NUHazV97qBybtPRmsZ
4ekyxWvNA973kIENQawJ9u8PO9UXHWtZmyMmtyec5Jh+iJKPkxVuaN4A4X/FVsDlHqMspn6xgI8Z
0mN8uzokdeMfYQOcqx2GdX2WmXyBZmuEvtImyKHyCgoqmdrZLmyh9VJQ23S5TUbd0bhB406oue6D
75XOHCTbdaoLZ5qA6Mt6XSmNtOqJNDyaFUAxH4G5pPowkbT4C7IVhcYVn5dp57SoogipvWHcvN1G
T9c4T4fiuMCCFp9dsEkYexC0Kauco5OXR3wyGKu0p6SEDJMfBBEeUlbLaNndB4HBtB0u15SQ2OVT
5j1MiA/vmvF/lqRLGONDYugttrkX+5WcOz/Rb1xY1qkrH/rSPPO8mC5oOdcIVzJWTwo5f70Ck0tw
lh/WRgndgybs0Effzm814pxsUEzOUzcZqUPA0tx0yowplbjhknVAc6UGsiSEtVs008hLeUkmOBXe
rev0HIol7UeMNBjR665JVSj5cu00zQ42cARsUf9yKZ3sIL1SMQF4OPX5POcQoAYyUT18ANzl+QLm
IUYrAEXUzY33+TcrlQ9g6gjHqxSWz448p0MLd5gfU5ATfg4LQ/HhSPLy11b9uA/ppP7//5EbB1vT
aUP6XdV0pQqomYs9o1M0/VgyIp0LyT93dglWwFLE+2Dd6B9Foj7uU4LcLyaPvGXtkxYTqQRowsUK
+dr/l8B2Gu5QToXuBvJzBzZKslcxPRkn4ywlFUWj+CzqfDrCxc+/wJT5cX+ZpCZ5s09N4RD9mgwK
pQNn+oPD72Pe3M0VDvPvQrnpjjgwfbfpIr7j9/pWBA6MdliCcRJdD6QZOTw9D6lHdhANNmtivk8x
qg+5DQSaFVm8rR6TnRowJhIAKbzghWq7jJ/Z5iAgKG5cNmkt0h7ugTZMwpmqJQLmcx8DhWbwV+aV
O3gcZxASppLI8tT7MyWcji8eZSuDDzJnjp5IzDF6g6GnET5Bef0nB4jHMs93Rt5MyFlipBuzqaOy
+bFUZM+ZpRTgYTls+0slAoSj1JSJsY+Rm+5D3Tebr60JsLxrWzw9Qn7o//clsqc7/1OJofg61H0/
nk/ZJFVhXUspkx/KSVTGijQJd/JjzFn3XOqZ+ft1E//zANhNieNGcCcrV9ggIAr5AzTATZ0krW9L
PaxTP4q6WGUlq3uymjIEIbX+aAeTLMuEXpN6G/ORr0Rjm4PbCDNe3B/eG9UTiARSTY4Y+pEdkolR
+ejl8ZpOAmCToXlAPbHWhhzX8BRlHa91wgrXivWmEosk2BWUNIM7MDE+WZEYr29YHbZrL+3XTScw
ylbzcdF2Dq5APm5/JjwBVBraDPjr+5sH1W5xMkX/dWmWoM5o7D/4fDjbY/AndPHZD3tNAC0LjeKO
1YBF0tIvHVzyDKnF+fUShyABmsVh3be+V2gQMA7IqsdZDUkQg8v5m7AWbwjdt+kqyaFG/BswnD0S
jbnE3PjHZvjKRX9S1mVa45B518nXce3AY/v83H+auEcOWmubnEADqeNi6wRXQNMUhdRvbGPGksUz
mh/ePPlM5SOoSNuLzFwd/dYafH95GYahNsHt9fQXgEW4+cFByJwgqOuYDu27Reg7EjT3v4RKcz6C
FLwPKfekV7CiZX8eW3kjxNdz/E3rpjlnvSHHgvFfGgSlqhqim3euWIUjJhTZOnv1GDsn8MKTEKKt
nMoH6s2nXCoNAtNVRmP+R5TbuJNPbJ7M8K7L0aE/nFuizpZC+rfH8PflXEFF8yMgsY5LGIRtL2lD
pap8qd5srvTGJssona2sxttpQJO8bUO+15Xtt0zoaPs00fB9JPBCunycmzVliqETYLu2DUsAdfnu
yBNit2A/RQA6thOdhjKBEX3lMiia9ZeHVtDWJJq/5p2BVkzOnJ5ja1IGkQgoCdxVqe31jWlXlvxv
XEUdQDPCj5g+vcJgbzGQaD6R5YIeILp9hG//IJdpXddxUPbH/RDzQX3JGZXIhgDlA8WtuPribkBo
B4ndV4uPjAXQYk0rxU7blPHn20Hjwy/PFNuqxH1ncslRfX7pwJNE1tx0ggOtU+FvuA4R7rodRGPF
2j6fK9JvVd7US5T6dgZifkRGyxVLdcHKfnwl/NZNUBUfGdU3c1D9nlDQXEnOrhYIzHZ6Vnbv31Rq
2sCwsHeJi6QWyBtTrfC+7JGNoctQwSh/LneCQHSABf6jxDC8tTh/08bd0fUsVli6laCxoqpdW7DR
7hiaNF4oEKz3kPbCNQ0XNPU+yotLSYSKvgxJKhk76NCWVyxx+CQ1fbfHJubhJlubrZgc6L4FNuYs
7LUFsmJ4eFIQKI67Ze48EdXmOdz2QyMSgOfP1usdNYHveKE6sq9CRSP5coVBmwoAGJACxqPVtK7W
Y6kZZscK+DDKmsMbGFPm23zucStWUFRN+RywTt8Qfix/haSxay6iJlmlgcxr941ymjPSxi1k0Kvf
u2ZuNVXdtilA4rc+NrCZC5xyuNWa6e1eX/A7Y0pc/OtmnLeFUB1Gu+S19wqI+98rk/lCzNg6XrB3
gwBrxLyfSoqzWgE2V2hqncmHQH6LttnU6hjL8YRYWeEDK86MjBs7OXxEl66rWGTfAswY8P6xLj/w
CHXxpMTRNNjERCtJ2fjFvMju1B07u8oBq3UCN5r/C8+YJePM2Uvl0kQL9K0r3+BBvZNp/xZ/T6Jn
eSP76/s5R/wi8Xw++6BXwVPdLfH9+ue3jobG86FTSWPxK2BajPkDK7OUkv3ELsTUm4r8GBmZju2l
A8mXWp+cQSlnTbjDOdDoOk0VcED2JNXp+GtBuVNycTpKpS/0SVp+qavbu7sH4vb9lmIA1NruNvWe
KqLNkvOipaY3ATdhundcQgYyEfoLia4kpFNJ/k43dpbv5Z+18Wg59vdga4Qs5hH1kxrrdvuTMINb
smDM8rSSRk3j/fW8cZOHa2qkc+kUJ4xptEnTrXN0uxW1pWJp7h8z1s+5+E9LS5LGraWCt4o4kOwZ
M5YCeyCrE/M3HTPnGBsEdIG9CyqMj1s333n7Fy3tx8h3l7HhxCY+hJNOnanqd7SUBo4m+mtlubzH
sHHCfaa1lQlX4Wqtp78UOoN1v+AM1hHQTsv4cwy5PCkJH+dtyhEEse88x6bMWAWT7DmzKZd7la1Z
12zoQpRv9FYCIbr/0GQKOUHb58SaXT0fQ5Ko57hLWvEX1ZKV5r45khsk7zEHsSlqLQq7LJMUKc/V
OTenGLr1Y/o5NefCFriVuetIX9SWnix47fZkwWJ/Y3tWeBtHr6h05+ApAXQmdMRsAc75HJeUQw9z
DCDerph48oDa4Gud616958FQiv9m1yy3ErqnfQ9bLZ5XNlBwx6umKwvVGQFnX5/te9UFd3/nOf2E
oBphPa7u/CEDLvL4eut11syAF0mwrzh6qSxLnThDr1fbFrryMjzwSPK3w7WUBtM+famzj9uz/xdE
MhclyNyse0mb+/9G8TxfmATAQstoZJ1Z822HXnaN6VP8rngKcBIksPDkLhQlVG5qlCQQaHkUTn3t
p/UYvG7EJLve5LZ3RbY0oFft551w+zVzxM7OmDIwhK2GUqzT8OiAm2Ln7a9KUHLENg06LMZuMC0I
nnMpXW95UHmQfPxY4o/D7l7IRPrEQG6K72pkc/E/pA7bEBLbEYqHoXksBHzT9d/OiBQejTgsXiUQ
Sif2w4VdvbYYjT73D8j7QaLMKq6/7TAnjAavf/QSdLMRJVLyBuGtG28SmFcdwieSMIvTbLDdotYf
5WNJilGsVxU32STJ79dttX7Y0fIlWmAh2+FS/cd2gcU4NQWl3cIYEe2vbPzo3DDflNx7BI/dCH1J
OFsEtTgl+nYAWpZ3mI0kdPDSMQAAZgsvmbZg9g9BLwdd1ghUWvu4dCYSq1e3fCdHja2Aq3USxCjj
W3h64XA4Yd5iYqQffIngbp8OpzLdcXF3HZbmM0mLbMK2On1G+9NRIgJ1Ya6TH+z2IbCeevOh9Iey
427XCjsj0gjXVkEqBYkkbD7bckCQJNmMW79EQtThoxlTbbgF9+j4IXj56sNhEeu4YDcxGcoH1m0s
sGfdRHDM9vavMBW5/RU7yfopK8ZluLBVEZSnB+4rdId4DETi1g4AEWmZRlTFF3tkQSBxvA7GwCtm
WH3XeZQgHPKE4g69yvXlsWTGnCLEac3oipGhsgRjsTU7sVbZoOPhW5W/RSaFRbj5ehpgXuFOV4WT
V6AEcIOwbk1fCFtltQjk7VhhtzTRz/8MwlyRiJd8W5W232fIz3qIzsn2rAxA4P8KOuezAZgGcJ1w
yuvq1yjYSkvb87Ke/OP0JyDkx5Iu7Zp/SzfTVSkLR+UgLo2UdbLIskREFohkffs2As50CtjDj1qp
7Rk+BfBhcUjP+Mvq5DWARTrp9zlHOhOHM2VW/xstFM5wxUusMvnlHLFN9WmjNRb1p7jfGyRrTSUK
OvimRSzhwQIUs1o3+fHJDcC0Y1LogG8TSC122FguywTooOgOkIz6vMxW0buHDzGXkO1I8fQAGHfs
3nhsKBMOU3b/9y5tDRQATLiNEBN6kUiOZKem6Tf4ZbfEUV1SKnbRwXjxiCd0gZnnS/vvxJB2UsI0
FKwxkVE6O6+fvH8CR7IhiTbIO/ao4oWElyBBVvRKZHaLX61SZeUpXK6X/l+9YRAEIS3uEuXMnIa1
gozA8d7Zzj3qQfONaX/L089YTNkb5O0JIzet6fz6WT9jT5ssRe2pjybE+IY1qbOJVEQ8wf/KWw8F
p/SR+QobL4dsQCeQqYLBoNTHzkOFFd+XAv3e6T6lG+EfemP2UgJgNcAU5vnpjVjJDmDsmA0YQesH
r9dJy/5TvpLC64dlJ5ARzvqQ0WoUr7KWjtHlpT9mWUJDL6+a0FQczd8Xh4cXSYc6c7NFva3c2RRb
81Ejyn1g0mg/wo4FoS3uRegC0GcBxmYorBO0Y4iD5D4h6PzgtTQkAc6o31YEOup/N2JrLaZIQzc2
Ln5Lg8RlNyS/n8gjGgzje+WYMUP0ILfSFWjmF+Q0sLdY8wYVutT6n6fdqy8+p8Lb5wCR86LB9vwR
hDltJDenotHaobJT+b6LGt9ZbEYsfDFMD0OrtbtP0Cj5TEKP5g7lL4Uc8jyqhlMN/BVdKOp8t+1I
D4zO/RY7SVWKh2oPidQ4X9dNRylx9Gx4P6N5vrYG+UxDITicwMwMN444c2aFC0/oEl2qROP9znJt
pmc+8tlO31qDyj80RBaksh8jA0y+n/EZN4zzzEjGnpZ3X9CgBD2dM5spy3q5YBVFJLyeR/QFrQRp
PYxALFoRzlBEOtLy5w6/2whX7LbgPTUxzYjl+g4p7GT2VojHH1NGyyR02V3Q3F3K10B60OUVLFer
UlrN4Gm6wStZiguvn5CgOjlRJvfSAr9X+8DIZHwYGaxykzUNMTCihjPgMrFmU7Cc5Wj6GtRzGUf7
dwZLyF+rFVv47q9zmT3Yodf+kRlVKJeG02jEm6h2yYCRDNOWmbj+mQqW20IAhVfr+OfVeRlSLp3V
qU1QxSXrN1Y+TUDG4RPD0NtOk8rE284qhLFxJbi+Gi1WxiJ8DO9umnSag0cbr9fijfLHORYdskft
ZqHGN4CiS9OpASVEve5yvsOU3yBwyMDmo2HCQCfYKF2sriNImeugOsXiJLovomiaq6lumMp5e4Tq
MJn+l9EwpreBTaHwWVm/AUHEm4eQI6fXB+zSHi9SYb7LTUQbEAcbwfcspiVRURuyE0esfgKnzFfm
TOaCznRC29ygm3dWfNCBTUScSzENuIxMWU3GPOystOqid7+Yfo9EU5lDH+R1HT3WnDYIhUCXNOzd
RDB0kJXsCeDyfxVBKFpzQTRxwZeGFEaB5jhS5y2k00YUapwlJoEsCTlQglpGP8PfR9oFtup7W7C2
DPrraFEjVUV7pyIuoLpKeyvNqlQuZS7OVUDDUuNnL+YniI+qCqvmUmctPj6bqc5FXwrDInhgt+V6
qCe6rCKnjLA5ZwLNFezT9fCEOuKaGrCfeSI8NQMQzloHSBB+kFjb72SSUKmF0NXbytBGp5s1FJOM
K5ehzaU0g+ccLULM7DQgiymhiQWiZPZZ4mjGQT04J6CS2kFnt/qYk2jbjxNYVwToWHIl0o8tJDOZ
Cay21iUlf1xjcBJx4XEjfZS0uhGwVoqlmCx1abRN329/it0bVyOqRpdcEV+v3+NHf6bXSlCHLUH3
8JaqTV2th+dEOoVXZmwTKSM7JCpD1cbMovEWdh1ANtP+NIld0K0WtRpj0CKiOly2v1z2pqkO1yEK
rkaElsViwvf5aivPo9HVViixKbXCIAjvifcsjHpX5jCNab5bqoTVMa3zqRkeaW09irmnUwJBSwo4
uzLEoadheWJXmd5tH3myWBa4C51gw/xnNtZ9mCeTbdw6dfuyB6iG7dCoz+A1hNN5+HdfTlr39CBE
qXPEh+Gc+FDcujFn3doLNNmZzKqyehK8M5Alny2E9kk39NPNm23J+eEKjfq01xM6QXC4o56PW5CT
eYDXt2zGg0nUqVDg3qNeNo7oAAzSkON379Sc5YMuJcoWYfz64tEPbBcnL+aeXbmLPMmYwyb5WJkx
nNDboFeWBlw9+13JESwP/veeD9UinXl5EADMTI7izze0iH9aT9eshOQDs6FmWqHgnmcVHJgvaf4R
XOGUUziSa/GbWbQknQ4XDtMD184HzXX3ymcoHDDA0tdacXhTNfqqIgA0OZZlQYkQ4T2Dted5tTqQ
+POVih2wW9wWT1t6ZharlTXSfsjVynI60Am1V2sDt8eHPBWKrVXa0/5OGZc+e3zdstX8iIm5+Ygf
HbZsaj/6yk2Z5v8lHwn1yiGa5uLyGfDiwFXwDVzB1pQTFhqgl73kyMIPd7owZr3UreJsqB5XAD7y
soWeJCROAFwO55jCoQPgi07nRmBJ+mUL+9DR9ku8bqo0htgMy+lEWT5NiARfh3UuUPzZ47g4PXcT
A3q3Xxv/vCmmUun+7qiglLaXpRIxM8DxkorLVjnr0pQwHhZILQpBOeD375ghaMQAg5gl003vkhAD
iaVDR7JQAIPB7CcumxGRSfbM/0D9AFWz65IzokCVylVjGM0BDJc1B+0lEHjbQpXZ4zV3SFZd+3ph
XOorry/kY3YzldPNA0EIDMZnpgsLsTplVghcoeBUaX/xxpqaXm72kxy/nZGCjyalyyHdrZ25WHm8
t2DuGwH+FI7qLI9y1nJ65jWoc6sdIEZG+lDFM8VE790+kc/xyS89z+CioVVEakHo/8GdB6byuFnT
0LmvBbqoHBI87YS/pUWir4UgOvEbS/HSs8efO0Ioln8UcunrUk3KLs+MJTUo4NJw9GeTCtelZlc8
yV3tVGH5y89ZNnOZayVqcKL2ghS5DJeNu3qWPBQkkh54iOIz5wr5QR9ruo4WtI1xOFYQVgDmLAfw
o1hU6aMSKK7L5HYurnwd62S8S6zTDkro/HcPJG0nx/8I301qOCAXmXlQLceavyMX6VNi0/2rpRk6
lpCGtXcczZJKVPvjE1e0ERGkEwpDxdTfdH9KmtTou12opb+v6h4L7lVP0kpy+VKftSFaQPUImqPQ
ESCq7yl3o8N2IsPluz0lbWRhIoVJlDfc++nqxZZM48MdnKVWXGurV6DWh8WJ2R74xn3cxdrMsq6g
rx/il8D8D55zLBCEbAOBFmcwkRlxOlsGy2YBbmiCzH47vHMk70Cg5ISfrtfawhsoTQGvJQMwZXVF
XMdO8iMiqe9cJN4d/IIiuRtiqiXr6OCqPD9XHtfvGm7wndWm7MgLsWS5P2/htk+rqmUR2/Vlxvwa
Hu5437inEKS9jliuWpslBXhd/UUqQf3RlCZAwH9Npz4mIG1KelS0nRaL26g0v5uRf137ZfGwujgu
YuuuDi5jqtcg38/q835RJPdRwrmqoYFZHxmC8Zl6/0/HCRZhtsWCNEzmg8TTzexq9azbvQP5q0WN
DKoIi8/Dxi/eqhksdhjnAO+NatgZ4fdxJip5fiVvn15bwNzEq62yL/IRnChOfcuDNzuPYns0zEgz
4CqCsdefvyYyi2+16s0JRY9nDOTat/fFO7hpjp5DMooeZZEfDw2eSGlrQ6bNOlhno15+DtzjIEgF
YirdQs2iCuAra+bKpgr5CnlIbuiSIsN0d2+V+anlBZ6EDu30cmeoTMl3cNxEtf05U4/vYjJqGF7O
3Evgg/v6e9aJFN3ABvEIk2iKcBX0Ini51q5ZiGcufjzb1Ko7q5wnLxJGxLX9V/y3dW2h3MQne6u8
IFtyCD1otR17vWtMXh+mmXg8Jb5fFD87i4arOOadGxu+SuSwvugFMOHFs5tlu1iCIvY/BZV9v4H3
W49ADi1XWT4hy0XsTlC9fJTb70vTdC8qcvQwEfSVYndnz/j5vuQIdw+mlbLMizTQllbzTQp+BrLz
h3MUG+oOWDza/QMgWzipJKQMLZD0CujlOTzC1L7bwxdK64XxEqoL+PEhMYbeJViFzWbykbHpC56Y
Tk5XVu9gaQjO9TkXyubJjUQSiJN8zaIVB6gYn6I8w2YgvXcSZtZv7A4HeAU9uwR+VFZaR7wtQgGJ
CxwiL1PZ3veB9EEFuo0P/Agy5SbFNmana4IevK1+QeQ49OK5FCDtpjzb+dUrcMRy3hVj0Eb+gkXc
Oz14iDOH0IgNae3f+l2gwsSqRELXWW7IdUWs7aeAZWrSzRSLHYqLI8SJ6WwbhaUsRttFaEpZxggZ
j5yIx4uFR9ipsi3as2bydJ/hgj344sLvfO3vfANyB1AcjRh+nbTZJVhBYqwSIzgvKytctCblMa76
4Jq88DpCc28uddDat9tfCo7R3Sphp5uc5jyYrPQUgcGcapl5LpKTjo6pR7HoI56AVCmhe5IRAF/C
0ZzRRQJRfTTFACOfSMg/oCCuX5RUgKNBkBf6Jv+oFKLGsHjoPMWvEWnP3PpeWZ7GEsqvi0WQGsn7
36zmYkzSyGWy3Dywm/rBkNZA/Gtxrnws8Q4Y7rc5jtqWH4wmIQKruhlpmccpex2JBA/rjRUHO2FH
mTT1gfUfq/URc+AJFn1/3WCmAvTtTo77drkmsyAQviWCI9WSIC7iEeg5Ns0l70NkWjWmscnXyIZH
gB16P9VyKdAgY20psFogccLakSe0A1sMcn5K5uLGT+srTFjhuZZd+D2D2Y8x3m7yomV0af4PvdLc
8jVDp9/3IVoWL5jofxHtVMuceCKjnP5Fxm0nKR9UHrrN6/0QXle5P+AneYHe8rEFD2ipyXf4oWAp
HvR7SGVtw23Dhq/9yLBEXvhQ2PmxusV3xZ5v7eWqZbka8V3UIl5lfBDDoySF5vdRBrWcUnh8A2Wg
YGcz0oZt4TxwbV4R6fgDEVEaSSgpuiiRSwVX3azvwiyUh1JLWjSoaxnsqOQ/QCVoLpuojvv4PUdL
e/qzLZWIkuAViPfD/W7zn+qUhsr8UiBvhVTLBT5aKNxnVBmDjLpa+0XORP2phvw72l75PZ2Tgpaz
scGIW/qlIKCnoEMaxVpCtNrkQdm+sfUx3UC5TvFGEcEaALn5fM1/FBRRafpWrJ40L5lhV004wssc
uzrMpcMlzYQwfflZi8iI51sx+FhEkqsZGKw/YansemmwlXTXg7AXEcE6m5G9YUOB5+DeggaKJao4
6JyArzFXJrrAphu85AVgAK1SkT7fLj3AHpQ8HRM24ETijRfd1culf3AKWE1VvjYDuHDrqISmELAo
aOtgwlpf++Q+MFt4WQBD2EpWeO2cIPslSH1n54gSCfb3xIOhgAmck43/fgbvq2zb51U8LZlJ/Ay8
gri90DWhnhIcQI2GQiz+wP63cnu45D0C8yqTIDQsYWyJpv4QUmU1/5RIXlIX+FYSE3lnIaRma6hf
+sf7kNgpY8Y1bUeSPBDrwZwMmU9L0VmwbGPGIaQa6TA3H0MhGtOc8cJccJ1hWdj8RKg6tWnLlVs4
RdrIfBMniD4YCI14yODy8ryqfvktWqMpLxPlmDbQA2ewRxc4U5HZyAfDkXVZIpUMedrYsZkdI7VO
sDk+ny6PkkyVxI2vzu3cmNz/GdEJQQv9qNfCv+EaIzLIg4SxUFVMe3k+xsVHzxxcSWz6r6WH2hfL
9/fiJRBnW/nTXey4y/rNFeRVNca927XxR3WlfXCfiE++8W4kgRenYaST+Z5z8bWdjVOUXpUtovhi
HDYwRcPLAPP3LX01eGWxmJQh/H1Iam3CZp9ws6aZ48w6st9fH0aRzjqmI1D3m0Wjbru1tm+S8Szi
BkkR1Mv4mZ0Pxof36/E3P14E8XojNR7DesN+sai6iN4sL65vu6AS2iDo1LeDNRUc3nRefag0qviH
RbwF6pjezncWu3gdIa3/l4h1gkXcZCGOTl2Zqq6o9wRcz+o/IQS2zpO6oMmuKu7NOpK8KLKNXXB4
nKc4FDht3QPABIWmA283h831pRA3Sy9xcplubYW2woh10R48vd6zkL2njv+4ZTtL1iPQs25RTpEJ
0z2brTU/kb3y/AdK84Zag1E5wuma9uUKrcGncyAYotl80SCQ+wZn4RhwHRmKcURqzM/WgA6wmXa7
RyruXOnJHU59YbeK3AQq/TJZeAg9J8WwNsVxJqGQHjGU4LgChmXa0ykORxezk6lU0eZ5qmkfB4Gv
pwlXa4dRH+LIXBG6o8DrdW8AOi39J3fyqsSt+504tG3smcE7T/WD40J7H6Zg9eI4i99eyPZcAyfW
h6izXRyQ3/Ie/RGZvwXD9ALjmpM/WcGocB/gNtfOCJOw7RVKXRYkGydgsgLYtvbcUPzzQG781GP4
B7ccgUtKv5bi/1T/kh4MumIx1+jNLNpt9x0aWAqDFNRaMB5Z0hPDrq2BY+YfRGBTrCi/7OsExWhT
DKVn4UdEVDyQJdSMIsTF3nOeXOo3X54VKlmp+4aDpKOIYY5+XapUaZd94iwl8pEFcWlp7eLX2iZq
aGnTpW+mk0QK31QpsxgFg6EvM2425Kk5FrWGlt/FwW1+LmQ1HBaJ29e2Fv7iO4mXwTkls3jxHnYA
0P077Xip4VgxsUoLNeG1ZE8bONAwJOIvAF4CbgOF7cLUrUChje2mK3AUBTcNCmUx48afy+YR6RE3
Sdtdj1LsTr6HKJWT0mj+yGuMYETef1i7gMJ8m9M6uXJJe917BYcG6J2JxdWQBBRc3KojR6ljwod9
zL+gjEDojJAVsSxLUNGBLRLY7+MVJ7fNvNVSYAvMoKypxkckiapPjY6lagmFa/ZYVuvyesQC859S
Oduvxu3x4GoDefXb+3xubEsMDEKiWvAV6wGphjeLBBaOFilyN0xT0gSXc1IRrvT7KTJQkD/3YmyZ
Bd120h3zYKtjbTou9fElo7I4a9GlPMNeHlHz/JXfZnbCeqSRzODOVJDcBK3z6OKVRkWzyUZIoSer
SmDsjNJMDP2sRjw+NHZeOEi0V1jHEoQL75fBOzcnY92vV5Oh8YMhuJWmrvqqWmvtEIJRA567Ioox
A+Vab23h6MPMTpcp76HMSzlrzf8O21o7ctvQldlm6YYLRjVJI8pPTi/5riUryWU6F/Gl4C5HC+74
XH0gTk7gFTZYi+kMskWdCi3BxWFrLMTrxdKIDc5dDJg0IjYmcapH6ZJY2cJ79/7NkTsobmcP6Erp
QTgraINj+EEqiCqvC6XiQ3unzDmNBbP7Y0PcXKrplB0dl94OjAtfvwg8VZTS6V5yBi9FeNymalIy
EyZU9CBdjThfjZb5crELQzZGuTzYp1/EM1yt5yJd2BkqcX2lZ5bChd/YixXcUcmFzyL8Bn1v9xYk
emQ4RZMJG0RoyulcNNmw2vtPvqnC/yIwFZYqpPDD7VQZ56TLZ3VGzPxRpIe4duTu5IFUqrcDGkxT
k/D5t1VRu1jRkjzkdPPAutoDFV9sFxjZ4UtxQxsrvX0P58d4PiJ5h8WelnqyoHV/QHN4R1tJv2pI
I35ioyc1wCggjPC/mIxVab3tL7cOKgMhPp5UvryHl37q7Kkuw3XxP8bGAAoni18hv75HZ0xFiaCf
6yNBf5AjEmp73xk61uciTGKFo4TTbcqSx46mzne9H6hX5cC8p4zcqBw5jLFO4gxdMExXIL7Q5Ak7
OVoD9+y6g1s8nhL9CKwvQP0IkN5WuV2Jxy3GYPdxvOFtNYgkBfWIQwFM8Tq746SwMfjgwZfSBbsc
P6pkYUQ6M5ohdMXTh8bJzmkG3sE93MCmr+5qK+PBbIXBbh/8ixc9i9hHK/Qm/zq3jTjnYx3x7C+Y
0MjkXZL49JPMvaXzVZK1U15EmjQQlIeyxHc3YzcIJyRlhR1PJ88MbZ0qW0foHYNlOu+0bSfpmfsN
87TB4GGba/xR0CRDodyag6r1PsTFy59eu4dennc0uejPbTOaL0Hm7WQ5mzok1bkbY9WQzs5J4zIz
wR+/R2XWXJEo4fok2yooTn50xDT6EpaBH8GtOKJCY+EWKFlkNkCpFdMn+BzVPMdRq9a7ZpN8wqaj
Ugi1l59xzixKwtLno3fbv3bIXkgWQ8uG6QvXaLfkIHaBJru/rIex7idu8oOmKuqvRsJ94/Sggz0K
OaoeFwNxnUVy9pGaiJXz7laXmA/G9+wn4LvVWcWvC2FQ5KIzhPdbQgO/ZCrxqr2yJGH64k8GE4ka
m1fT8NG5BJ9BJTR9a/YuU1J8krLaNHzwni7qBQlFxpfWP/So2u5kFrggpOBVARV+OiLkRKIRm4V1
lmMDjqziai4LyAIi7e64sP/jPOfnuE+zwTpvQYYaYCTABmB/8PQzoRpCi8ej4RuDLAKUuzSA9dhj
/XY+0YK+XxqNlvq4bx7jXjg6UceerJisZrBtXsTn0kX82kDw23taEQ3u8jI3gO4InoFJhpGTts8u
8wNonVR4OjPYO2LBK5H0bD089qmbP8LtACoWnLdAZDQrRZkMM0UoPLysAYi4MmHQzrFQgA8QKGGf
VGxRMhtPXx6thU63O/YXWvcmZiBmhxvnl/XnFu0Zkqv3YaXqU/bgjbRCZOTdLX/E5wMrH5N2Y9jw
rn0YM8dZy9tTxQpcv682f5huN61B5k6Q+RDOsLr1yGoQU6sosFOaXLlQCeuFQVbr2twyalK/YQBX
JLyf8WoYK6XHYMe3y+y9Ha56dVIx+hdvBUT6dx7/LKqztKan98CATlPhTojx4xTId1AuzH2hrCV7
awlqM/a8mnlP2PupK1GizXSMww9KtEaw+vnmgcCWlC0NAFxb+B33hCmAtCCO5M9qDwSKA7axoej0
5zMcoyg8Aj9YOn7JppZ01nYG8/Z1b3eceRbTqQ5AvMc95yBVyywJX80vrc0UiSIjfi5mS44Y2WeM
vD6YMPbHQjaMIe1hZyZqS+CAQcYWvZe3vNU3CuPtlBDLw1hiSyqG+Mli2n40FkzvQKDNie/R2P4n
+qthuMAqbv9d6XcnurZAFgXyMZrKujTxAmvnoKJnBv1TpkyxOYVkT24NTR78xxRFJmXT0B/dGtSn
5ijU5Ndz8VgP5Ng7FR8Couml3Kdkr1KzbWitCHJW0ylc3gG6j/9G5+r9d21N1QPNn9RPHmFW84WO
K1fkxL9JoSpwOfOqeG6Ww8xHge5rlSMuGmziKkssNiWgO0AlXs+SkjlZI+uYfXhu7Yt0GQUSnOa/
bOZFjIhWe8KGmZhYdD09eyY3XIzgzURPdgxYNyzCCM0Ftki1HxTRd5oMhTS2e13KtoEqq7NJTtZV
KGBvKYN2SEi96I6k28/+xhxsF9oubrGgNIqIB9NAC5JVcfvljMFunZCdMt5iM5By8Jxc/BZMDOX2
3fOd5WTFkgUH5R7GSB7BAmTwQ6ddAfdHONfhcFG8cBqd9mJ7D1SmUzlCZiGYHgtg6PBjk8MYRf7P
w3imblInUF8XnDflIkHpLSBLvQcLqeB2Jpx7Jva2TxWTEJBm3OWEfM9ZBNAfqwNNn5WKVaeqGxMW
rmehaRHfle1e1v9YLXi6QygtR/B/EjN0hPT7akQcEXLgCQDWrq+itIqeejWfbAMWxru+Anq5Pkxv
sxBDh1kjos2xuPxt5beEqPAaanNnGS+qh22vXnxhLMCZwc1US6oyDiMDp6v3YQqCTAyTuesCHLv8
qaWqhOvbmyhvDha9JyLw9LGRWx6fvJEEZ7Upgck9W4eLlQXXq+z/CCiZYbJkEAkWCoHVpjjpB/Ep
DcdzwbedZwGTKf3r3DVOUCq5gBBSuntqnaPY/Tnn0RgySg9ZGtv9Sac1d2DjjXq5Ixa3RY+E6xkV
Wn1mnNp/fZCx+AlZS1OfAkSROIqAfkHdrsfuIymB/hN1b2JItsV6OSpbRl5A4WxzazxN/D6aXdtr
R+WLGRjctAtENfx4gMUw9wZD4z6I0jHmWIF9J5QTMN4q3rVe/Od7nm6yuXKdXAjlzpiewY619uhU
zSKQ/HL8monKRLcuPnTvwyBz0vMjwwxDQIQOHZVmGLABAQJZ+s9iD8++vipLj4ZhZixB6TNspYMH
sK1uPbL7tSzUPpuOEdKlb4m6uRtphtMhkLX1TPY+swSBXDY2tg1wDOoTg4Z0oZlGNShstVYMv9lc
amuQkUfJfBV2Uw89zbDhy1Cv5noI62tZzs98p3jrUdq+MpUqcQ9Fi8Doz+BLXUM8r13mbZGTLHKH
mENFfFqW4ip7tQY/h24NhY4gHFXp11G6C1kddXrJ1d8jSNxflPH6copqspNJNbiZRcfQnndUoA+M
1thPvsCStXnr0b/qjVBRLY8WLTvGViTicmyuN4jGXEjpdyZkQ4J3AWGcesIdP16etOVENcpUpHOp
6q8tfxehGPzq3Ows1voaRiOLZAUxSfMPBH0gGFPgdEWpC0xoIKmUkS/Y7/lZmfLVGMXaHd89RAGC
w383MtLuhwWckIQfk6evTof6m1qicVVEo5xQIAIQm4gHKQdZfTkJ8ZhXdlGFyGNQqy4HQ/0wSL1F
at6U3vlfcxUBTAc0CvSctiYhc5dd+fvdCzhp5p0d+MWEk+aj2RVYmWbtKaFmPr6ny77hLzZUT8+X
lHLpUDvAbkhctpVUDJtjGlCQLJqfJyjVS6zj5mZtYyOLXrxR7vAtYHJ076goe/+AYHBt0XgZLjCz
zklbtiAyn02GbeFpR4PyO1bVROVkDS1vpN31NIgO9+skH40dFsuHQr7U6diowzW8YyoXeFdZcQif
BPCNxOLcqdrnl/2oVygnHqFet7XUCOJZUW3CynURKoBukoNKrsKyOFPVbXU90n9OAd5X/QA9HpxR
wtzkwCQnAnuA2GcaXA2hvLdg6Yvm0TIIOPOMXra0N251IYoc1oG/JMYNd9VySyVrJh7MAXaWTheK
MFlOjFm9nq8RZeAxpykyBCSbEYf6O0cnkqxdxohxM8zDZ1PBlsyx4ZwEAulZwBlg3JuYPLbEugbJ
eRedWq0YNuwmj6yxuaDy1lu7y8VnENURWtBkJL0poPVBzuyEITaEHnUf99x7TL9eDp3coP9tFmMA
ezCc/SGsOT/bp2XxYu5d9f5QGz5q8udd04uTc0c6VXdscdeaMjHr+/WXZn16lE2tOPTulvHeLuqA
NVM/i+Xy8MzthdaGy3HSX3d8oYafQuVYISg/MgkPPBulpKYLE6zeQp31Eb19YG0pLHfPSS6onUGh
ci0iVH0bizCu+LJJ5ypFSqwoYlZnLaxqDXHzibmi0fMjgNiPj0CNjwgduwcKfr0eT/VyYusyTl4j
4d+kPUa+sgumx05Gs7Jck8oeGLak0dmtEe1WJsUpcIO09d+A/UDrj1YFQLnyXps+TeGlzkVofG21
AN0pkeHB8Hzaui9r8z195sXZUOphVdZ5yUqxBjB2QWNk2m633s6tRJomR5Iy2G7VL4lW/9+o1KTg
Yp2/z/7wgKXfLVZR2xOl9PHBWJkHkaK2R/Hi12p8a0xurpq2uSGf3dYZbNajB9yx7rArPPY7R+pX
8Wsxb4ppJh/HoEov96emY5d0D7/m92ctbzzMeKwFxfM3vUJBjnjbTKhCjCkoBDINn49gX8m/G/lK
RYwWXFrMYJFd3L9vf13aJyZqGwQE5342MzN8A/XNj88oN8EK1jLAzDJCf/4I7n6pdzMuXf2+orIc
nWiVESNtocDeiyMeORs7vYzIwC+1RDD3b19GgdYEipfh7cLg9ffdVI0aYymdrtKoEdLJR517iAL7
KQ2lvzTVvbiOwnxiZIe+LoQGkSu5NUlnFfk0xonUWSMO296p6HxyOHd76ZVwGwZ6PL5YsMpHRMfC
C9CvLNUPQbGiAdtISHGHbNpUT1uNXP/6ZAGxx+avduCw7A/+M78x285s/Y8oG0dbZ7wR26Un18RS
7IhthHY3nbFPbi6/4GNQaDzol1mXT0rkCxe50iso/qBz+OnkmDjfXVbsRiZOLspHQWKKVUQahsdw
yqM0QuKRPXOkgNRj3Qwk/v0L7aBGpYmKh08IJZPmUD2rVHfH+VWarsA/c8rpVYF9WCA3MQDTUa5k
SFk/zNE8maXNavXYMGKj+Itpy0h/SeHVqFvWFiwjd7altlBtezGnBflbHfoiSsZe90/MVsFCC1kH
2qhzjyaF3edP5SEvfewbSe51u7EHZzUkMlt0G+iBbwSssqpCS4zYgXHJve4+uK3lHrJrYaNsumm4
moNIrQPknk4P1pgGdo6qVFkgWkhKaJMq4KclcLB2CW6jovs1/Vle2ZNcZLlpGXaYCLthQyXv3qKA
kCLy6Movrsdpo3eJhOUxL5yiaRQhW/eYL9n6hFF5SCvqw4Uqp4sUl/Cuasv+RP7VT9i9yjnCuckd
V5fkwEJvPSjNdS+1uR/5jKvPtSMLHZUVR3H6Wi1B/PK1bRg0sTQEZLjm6qpGVbTaTE5cCfyeRClW
vvBKo/24wTa9RfswUYxI6U8I/bF/ybNEFqdJJlFZ0bp3DC/GL4BLIch4VYkSMw3T1/swZ03qoNsX
vNP4xv5ICRP6UJ46EuprPXoxDJIuf4FvnZbihTFPenpZvxRhky8rM+eSNANbuJ9hrQOfqgPjM2yc
M57O7wwBpQpQS7jP5bimm07ctaJBsATip5CfhuotrdwlDORCe+LEFk06xB2WtbySwm6uD5atFaOu
+jI2+8uPyLurcp9Kp7nJGw2BKu94m7KL3JCvH1pugMv8M8VPDO5pConnVUdxidOYlY9fUxldjX9A
vuJbP+xCgLrzwuR8grb3elmHcfKLv/9SOMpwF+Cof2SdSfBSdxKRL2Ccf4t4oxa95ProfXcaCS7s
sH1RiiQqE5YCM8U1SIbRHgWOEHbxbY2aVBWqL2PG5IlIfLoP+Hk0fPVxE2b6Yj0uAG2if+zG7aO0
WPK/8+ue6ZnmofGc7OThRzUWcaNlG+E6xL+OsA3LLzi0QBgvd8KuCasOgLUXiXn9kNv4GGXTfoE4
onX6JGuDuUoyz0CzUhIMuMAi796pyTTUYQz32IP/hkYx2uYrNprWr2i/1YWj2xDgqHtlbe/iS6ix
R40M2aeiPfHjXqWwcqLOqUfWNgq/nyRoay5kIZYd8F83KG9rMUr5AFHPQd1nhynQ0b7w7RXyJtkv
MU+HU8HTeHdULWCHeJmm2lYrDM18E2r64iMB7BvM20KXDJ+GzBKoKD3DtW89OpzLaDVCtalkOWH+
9dcWDWCaTP5Bld2wCmIX2pw4Ilb9pFE+9ASrty+DHRAsNvc9dXRXiUN82GnRRjMkPZRB0wWjbSVm
MP6yk1o5bBCGLfKD4NfHrxeTR8En1gB32hlyeysBBkmdSB6bqINdsi7wIF+UdZyIqnVU/M9P4+oF
NxxrTNw7ll5pY5EiDE5ygSrV9hTFRrxPiBFyvhFZdO9grMSQoDl1gw7trlQ6gDx8gHLJgXfkG2h7
XwuMEk3pPZfqJ8zJk76gwRVa7vc3kCPPtg4CdToeyT/9N4VMh2I+Zf3mYTA5aiZRim4EhWb658Hn
iCxzKIWNfeedaWxd15JrbaPcP9b+sYLM2V2UWzrhWpEgehdppQx52tnrcpHlEPY54/0UFAndMDQm
A3AkV2IqU+OhXnr5DQ9MR+M0CypqxOzHoN0nEjbdRQRuO5Zri/s8pr24owc4aQvnnND9F6AcCnPK
62AhDPvfYy3tST4X4voZawdYJmjqLRRooDhdPG+LkEIVD++29Q9C7JSjFbkQ1qtXNW/V8KWXA03O
jCbUoGtjuktbDyQ8m8JTbBCCuIwq7PAEyQf0HHulkelm+vmNc5SEnehIzLDJJnnoRwW1c0ZkdJxK
p7w3DV2CRVWSQC/11JCg+vK+UFGNP+ziGdY+d1Yu99fsGc0Rv2pHUiZpCqC9k/QM1q3Tma7UXZJ7
ejLVvI9jMsBJV879UQ1mX8GEs9bcjWhxDVOjNlnDl3m3c7CsX7sx/1ED//gBpJwCRPcuh6USNQqW
Fx/FPpw2GztUfjmrKin7sZxF9HDvMZmXzcsl5TOGOnrov/Z6Bi3t5SN7PhjTIb5MN45YWFXB2wKp
Syih+60lesUb0fVkhwLvoZx/1+9DcwylMsvij9cx6ZPrWLElzXzf2rl11Nq/GiuuaAa4RCXsL6eH
ElPo7TFlxDaPvS/aMuksDKDtMORWvwSKbGXlg2BxmUDd2cG54iPOVTEkgaBnOj/AjR/kc4Y72kT/
qVZMtwrH7MN4JR2I0rPH4Eik/ECM6caQn1ldunpokhPyLOxrPQwUkxgTI3JizysGKs+J+zpuFK7S
LuC3DLVePLm0K4vtt6qg6c16vc+3OWm9W7t4DUvFiPdtJRwH0oRea2yammCKN1S11pBiat0V+p/4
8Fnu7M1t9qdqvkk9Cr/eCy/MYl0I723I12pDPBDXH/boR+1JqfDVTTgPiY8Yzb/VhVxKygwJMZF3
ARWONP08Z5/ETmef41G59hluO4aoNVIpgu8kmszGT0rpJ1OlzunqPsuF5/uvuO5UyXHKv6Y99e6R
L+/fyiyT+gqK1vYYJXx3q42b5YcpEpPDfZUk0sDym61RhnGW6uCueHa7PxP68pCKXqMpYg+cboBF
4+DM7o9uQTYKGJ6je4EI6gxRhgTQiyHgVq5uAzXCd3DN5MOsiigMaaEQGd17RSOM7yt9xGPyogGS
oF/8xATJYxBraa2b7nr5myMR662bXW+cFnPbqAB+khlb1r6xao0zdirptrLDsqs5rJ5aDO8YiUth
QvDCDGmBJQN23itZWPF5ckBPD5k0V8e41zG//0btExP34lnXhKzaLfqVNxzHLo1UYk4Y77beModP
77cE4dAQlv9fBn+YN+CakfUVt2s8FPhoe2dE2YxsavZLkqAKyy7/5MExnb+YSy9w0q7nFxgEQP6y
ryZtedFsD1MgAQ6Fpgee0J4W3WkOqffT7TDOaIpyheZk4vS4kuyRaFFFu75C0iLCN/R8mztKEJAZ
y61povVP3yQMIKX+T2Qow0T1DSQwDgFs45moMDftxScP7pAvhDyS0Umz5nvhfFt/2f2A/tXhnE0x
r8P25fSEGcmIyx3bOaToPNkyvhFwk798m7wlz7oQujgzAwLByYRiA6xsCRJhz6ETIU6qkZfdVzN9
qXdJ3KSyRvFlRZxjCMz6nOJHQfg/wh0OtDXIsyXiUMHBD7K39kDZ97YVCOCTRzdDR06DbF9lPpF/
U6Zhz5zx0atZ0nm0bCZHnCCS3PYCkjOQigJh0DLCx4PPjP4RVg+gbGnjkR31c0qb7g5JvaxzTSMu
DhNx+ahK+ZBeG2HCZTfwtU8fmKUMXA9W+yyyft4QHW76v5UBPD+a3dKHLOk9G4xP3k8lMXS1dKvZ
b/kkwE35NHt8I9afWLEkhVbwEMHlqe75BP9lVsqxAIdeZPJHz7fRtz7LztzBhzOv4zXK1Fm760XD
Y9Oj1NfGrh2NpugqxHTla6iyzOpUMzjYs0fhIpDThm7AvW1FP4wKminRlMGjUFakCMRPWHHnjkMI
CxiYiQjzwUbr3HuOlkZGP528tnD/9J3Aq6hP/oqPmBspNRtSexGtqqTxVEd080IgKwXLBDJ3ChKj
Q0uOdaZrfjzQWrz8CULUr7rVBXoaSbQtkpBypeb2dSc6cF6aP7jg8JfwAATkq1xOwzb1BgeqgL33
Q0LpyaNEz9h4OrTAnPlOAC6RSX9f2EyIYGnaMBaz0wi0qGQckYVC04XCgql5WapRZHmNzyb1ezR8
XRBvkEk+GqtzqrfXYqhVRUi+CXmyddLd4JG3a+bOwg+Nz/dMxfu5MAGjce7ffjumnKl7FFC3YO/C
XA8jlFcH5nxHS9kGg4SqbyArpWhO2J1hu+XS0TQ0xtHhJ0xr05g0hUCR4x8UWYiM/1CkPd/vaSIG
EZccL+jcFW5+0lRzZIVeXfxSLNnwcbA6QciNbINiNWGowJ6COrlDi992xKXg7UWD901kPKjbQ3n5
DaOCcjwSHJDj3qzNe3bW/2UhxnI7ja5F4QsopvlL000w5OUQhSsRuBG7SJkrs6OWMyg1U0S5/59V
dLjv2R2BMYk7DO6XqUIZ3TdDEsri0OjE7AeRRDHRFgDfoHeEKSbRYzQ1o+qCgxgwwXBFTWp8eKGt
euETIrxUBVR63++qFcBDk3NoTqNPFvxBZrRNvRFmn5XBKW3l+O31nT/0tFr4z4jtSLg18554Gh+I
ptIQ9dpMW2i8CkKjdBaXbeglW4O/8QULx/zpxb79sJBRKiAA2HwyzOb6tVQ3uan0MQESzhjwDlsv
Px868AafaVMmo7MNkCwwWbF74dEv+cSBwg3ClVnL6Wc/bsZ82qyqoEzeCDwqM9UGhF8srlKamWKE
dUrobbQMSPIMM+8Ci714zrP6MLvePsJAbTH/ymsgc6L0GfB2+B2EXptkL/iiD+GowAsRlLSlwMHY
ReS7H4IHpc57UOPAEwijZ2kQ8VojOpyJU7ux/LRgjn9v0RwTFfKmj/u2y/+fJPCdgTLEiZBfFGK0
aM3aH4k3SfjlbvMrAW7az9+F8osKfNVSTBgbtVauQFmzcoeRRnv0cLx1YCb5WwdqbDO0hpZq4JGX
iDSACwgYV2MmPp3qBUYz9e7Ac/pP3L64wH6Nx6juoucRvq2snYHCLhk5K1pn5MXGa0spsBr5DkjK
V2N3TPd3FDOlYa4rYpisJfeFkNQ/JqVSwSqn22Xn7i3d2PdviCw+5pgW1exkPqCKgryQDquR1sLq
jDztz+wLDger08qSQ6RYUPVZ2u2yYIj8KPRs07NXm7qXc8jL0N1kOOB9IOaTMPom8MEdM88VquIA
AYDBwGuFwzh51cOhLPjPmviNYqY+eoIVBp6uUel/Rew0Lx5Z8CcOrzlQhDodm21HmHuLFpDA3rEU
XI9c0FOab9s/WTHiTB7VPFc78oH+A8QVgy3Z8A990wYFIB2C2nRPhCyvN8l719rvvBWoDlp8JMkR
FkDEaNf/QKH0aEjeHItYfs6N1002FQBMCtQlsV+LYwlTHHH9NpYtC47Duva0npBVnLDIm4hB392Q
i80evdLtQ6q5Hjgtie43mCN+nPFvFTlh0ORST62iDoxKOCZp5MUNdx4B+3eWCzZOya2GmlFW8RHn
Q+5PJLJyjwlse2XF5tkPO/Z5ywRukWIrUWyUaFE4SRpeZtijZZ5XJCdDgmkKFTmJ/2+5C95aC5uH
sl3Dlx6nxU6eOLid5I4l65QjnZBUEEk0PINYKoo5w9R4JhahOYbno/t6jdkTY9VO0qZyv6+poONf
R5F79nAuzy6Zu+/VBNsnVH1LN1aLsi6l2E6l0QS6LOScxyRsIDL18FmRVHR1K9SedYpazn1+cVO9
bNvw3KBLfCcHWgJ5lCAF5WYi6kTBTBh6u20wCBegES1IEwd3m9IGnoEIuKCONBYOPvCoALUZhQ7U
ZqFsIkdLd92oRxIrpXZgFW/FUbl5HGUCpzRLmE1PlLl1f4I7nsiLK4rNT4N9VREJPj6VCBNLGbHg
XYZMhhVlyNWcDpqnm3JRPUgO7NgweUta9eHabV2aZCNQ3yVfkwSsrIkBQXoNwwStxRLIzIQBSiDK
ejUpIt12AwKAs0zQlydpeVxospu8028Mn5CCAdNVdoK+lZIAVvjGtMB7fH8NZWUufx+AhU0zGmJD
Pwp8y9uyDaoycOPWRMXvAJ+AulpcefPbqUzUgjKzUdxj8X/Tku/WCO8ut7d2/gzSenW4z/5mqUj0
SQ2Ikv9MjN1Hc2piVVw7rb0q4NxmDe3LEddHYnMnF4qsvXj6n89w3nyA61oYk34e7JxgxL3lR7cB
9zsAbzdhQ1mgBeWNh/VSSjGkteT/Bpdjj0L8EBnH74rFnYekXGeXUJJbJybOlh12GCXwf/5DO1mv
GX/P5JQlT+y9pcbhymwnx8TbY1IfNueZwQoxYKXTawqCI1cNGwg79p9MPefuWInMlcUum0Hh5jay
NARHQqOucbcoFNvAV4FYO3kG5Cj73sbxD6e0gp7JyKCnUU/NPHSYe3TthHy3gLMBhyCfSlspS9g2
k4MmF6hobVgk6VCRNdEv14OHLVfE2XbKZUfn8p5sNYAUbyLaUbpIyxPY1u7i/zbM3S1pLp2Lturv
2fiBlbHuWTSe7II6gXqLekmM2SXzPE/xFnV1aUISCGVNeyULhBD0sfyEua3g+A7lEyF5D4qTjWYS
LW0RHWKcBn0CQ4J0GblSsXxKRUoQEXZzB4V55MjrfvrEwS0TMMfxGa6aO0BGXoRMqLd7G+5E7PPs
6wIGeEYqhuJhIXN11viwWozBIFF1UoO1uBQl1wbRfdX8ih7/OjHNQngJbWaYACMBPNtiXaQT1Qwm
osj8XR5kD98HyurkbUo2/YKErLWfL5x/6otBd5JO7vf47taJu01c38hn2R99mbV5XK8ejRLANVHs
7kL2DlgtZf25FItsvdNMtqcnnc6QnXdiABA+mvtcTb0Li3xnfZWBMkgdcZ6JV/4Cx87Jd1zzB33B
k0wwn2QB+o0aGOM0DvtM8BBO6DD4oIJL5WkP0u181smqHqeUYGVY2zscy5FyunFdvOnQdVECjOJ8
ieZZvd/6b3MToF5nYIcH/2IjaYiacONTjrUS+TCStgOssTr3MCLOK0TQNt3SmnjFQuzpxHEwL6uK
3Ql5UIqSA21hdtm+4J0Mpv87HhggEB2soaJlW1F+PZLQmW0uCFQl+AdD/Cb+H4o5RSPtM/valF7n
/v2BCrdYawfJ2cVS8n376GGU1ehGq9KGjqkeBfMOk/b2KUJehoImD+9hdOEUT14/gcOmIii66mSU
poy+17YgJ4bzO4UlXxptYcgHxSjfk4t39hcr8KrlV50YWT8n+U/eSKF4UosDY6dEzcMrKOoCcBGt
c16Pv8+CJrYg/dRblkNFW+xDb3sg8KE2a/NtyKwPDyOynG6JZWe8sGdmsXcVp9nvRG//dXpoHXeF
LgQnihs6ki7uILcbzfzxvXycF1wrD50cEwmJPIzCFY7otigwuqao03ElKljT8l+LMibO0QCsKEcy
LGOEA5NLGrZ/2XZTHqyy2Tyd95LRBtBbm9NdNyvccimqa6YDuOc05JvjiiuqiSrQkEiqqzQAuKdA
2YeoGFjrQrZNHnCWiJIf8REagqT9XBSILQn7DLhIAqsop+pwbS71VA5WhvRWESWt2wPvdAsdqxA0
TO5/9d/On/1e/rX/3qsAgvrYs5eCXE6Lls8evEJdT4jNKnbgIHQjDhpZ2eCY3gDRyOwExNnrI+tI
d7LqFAIYsoTgOEwMLiCHswNDCy25MfBsEseoIBkJSeM8cN5jxCMzvnLv1ET4zrYXuj3iGJXVo5Pp
GjIRzTzo+zUUhGLzLhM4lz8vhX50BBa3udlKKmDYpMjvqKBj8WPQi7QYAauwDUnuAnLPl1qFUBDi
8Gb0k+0UX03WHDJLxTItKwurydFHEMC4zBeObS862EIjQt8/u4l+QGNueK5hyy2+vRiMNevCOHFQ
Ft/N2u+VC4udajCcKiIqzFC3ac9THeHqZmu5kaMNZD3D8GyedD1zOW8LpQdwhCkGUsm/32TTmiXm
KfqwOtQpDt0a7nIfGJYorpYd8o4rTMj4fEG5RC/Igl9+Zuo0TVi0deXzDR8/aK5aA8/Lx6O8LMr6
xY9wTm8mbJncyawcLKqsshhDcMrRwWw07fgnJOAFUrX8x6CWWnFrPqItjrnNPQgyKEoWNQAORlXf
FU9ofXI2LwjmsE01Gma4i/eVlk01ZdYFiHOmfH/BEaL8DnxnQIR58Zooyb7QZ92rnZkWKDqwbXhT
TNphLTzK5aIcmeIs3R6Quww3mWdtuBV2yTQkAq4F5qqd+b7/X2RQD4M9khoL0xdPhOQ7dggkH+aG
fOw9HX7I/T6bWNlZKOCyNfphE5GncFDzO+S15rCkcz1TRbBYlXCo88s/2/oKty5CVdjgM6Oyje+W
pgC7PplI+5LpZV+YUFNr3Ex1thqiLTCXQTPvWkKfURcDP3OGcPSd5abNfX2Vyfc/td2C/hoSFZCK
Ys/SSeWogA+A5nE7WTHoLyvIrj1BYa7jhWZ/XEuNgCEasKeSqh3SroqyW9OKSMydUsmqIZRTUqdX
ZI4n+JgfkyR4ODE5E+yS6s8ExQssifchDvyvcSrQ49MwbJS6uIK5awEBCTeTtZ93AudoEQbRAzYa
S/l77OTLK+7lLEQhXNXOTmO8mXvVx//9rf1PhOYNwmSeBq0gOgPoXK2+efyWZhGAegjBMuhD2/Cb
9RrCMtPPsXn17O4Jyt9/ROvNzcXeeqF3U1rOuzU6lode/0QvPJlSG6OjJokGGaWHqGhOYfb6cy0A
MDFG7eSWGufgg3SW/UcQFLvSBHkpDtDUXucJ/XaKkmO+uQ/ozZ355tFahOmQVXZxhEHE0K+xtUt8
6F1P1wIYHCAnxDec4x8MwdWLCHIv1KESgM/mZUZmAfkieZ0/sM8Ln8KT6xq/CnvAqZkGQNh/1otV
f1u86QWuQy+aFakLOMs4QVPygiLyIgW5k7fOnJC5QiXjKPTP+vPfyNeRRPhqMCILyWFebPWvZAMo
PX/dotPa7BdE59WxEUlkUVgli2hKNYqxNu+fZRBxP77K7VuLThrOIG44xxgfWpvvz5h0DfJbVUVu
xFTWLXG11CmgcCnp/FZJ3R8ubcC4/dc7bXYGAI9ROh2D2pn4SOww6mv9Iit8GKNHbuoRLi3BGufS
Gwn0OGdNE7Yqc0dXu4OgQ5XqDdvf78qPb+a7XZ2UdMo/LLNH7g6tbCLlIJzDXsNeeT0JsYcw4Tx3
0/SyHqz59vUevSrdeYwViWruM+1UK5Wl9DPIWuCcoGhJplFwgwUcTVfP7pRnVT+S2mfpwo/BXUTp
jFjT11kPpzpf0nztwegWsls0kQMxFxqQ2UKfzFUpg/1G7aHrrWeAQ0WyKEX17ORmGntim34HjsEj
xC803Ro1VnqYmz0cux0iKQHKR+d9LVOLDqHBfcd8lK09PlkEbD+fjzphEqMQtzfLqHolVtCdsrqL
kSXLcIEKhl5OGFCMLjtj3pbyvxZkBqgXRS0XDgE0zvwtZCb3X7lP97yPRSmjR56dyL4Ed07Z6zwN
RIhKLHODtNwI0XAblhWjN/qE3HI7MPmaLGeB3Y5YayDbZzzgjbJYJYry111ZtFQHfx0xwO9yYEFz
m+nCAvabIu7TjMGsjhSqNTLzd6kIo5i5nC3+2EelCM496Ysh9qSj9jgJBYxekmRe/azgicoAXB0D
CDnyjvZS8u5BE1YiEbFgj0KgaDc1m2B/XGJV5a0h1h3XRWDPUYkHQ/1dzMFfhbxeZU5uUQApfdEb
csXOGi3LacBDoo6PlqVE69p2LVohT3w71OmyGuqVvWvX4sB4hECe3dSJ76IVNPdhG2iKWOs4bMoh
ztWZZHaA1PoPHL+CB4jTzyeWdiXpSKrkdkMEvd1YuVqdZ+zJYByW35EOSwY2eV7x1DQmdYzON66f
YhBuUmEFxn5BpcPTqEGSabB9Gwr08KDRHGnYnHIGAH7w/M1xnxAqNWswavcbAQJUk0NPT+Kgqbew
XXIwFVBMv1Vd3y2SRYNnCC7b4ZSyflaZNhXRU+vn7xO4YaQVFxmZmrBQ3NM77R1PKYXNCc/S/x5V
2o4iUrkjFnqSE7d8vNuuxjVp3U6b0cdUgFIrLocAEg/GiPr4C9x0oJiuheb3TRE27xX/jLyBmQpO
v54TNHXc1UZh1y3Pg8286EPN1sFlUdYK0trB7a3XG43sHevB1XbaZU+Sj4lqU2BMdPDgGKxiwcQX
30ewZFv+BboFDAyi8pmX8HZCZFNlR7OWfCy99Qow9HSIpbp+EioJhdz+b9R6Yj7R7aGKqSBlxYAj
raP9fpbDwM4DjEr31EuvBbBlRbZDPqap6otUX0j0PC1MiKYISqjUYfO03j2jh1XUhC3qFfvbhGSw
AsP9JVSs/l+g1i5SpGpQRDxza9D+hzAiYPX7L/M0Uvqx+sX3sxGfx6MTZytK4jOotdedMhgTsNhv
hnHls/QMccnLQIPlFNbzeAuLQQXy9Bxspw+9LKjoPE5HHqsxv2h05oVj+mehlBhmwHO2p7WCyIb8
4FcT3W82J79xs4qkye8StddMWV5UcCPKmr9FamwVz6aCEUAJNOJLnrp6xPgX3cn7zGqp6d9XPCY5
TZn3Q/2fkwbXnVfAMWyM8aNgF/+mKY77HTHhQNtz/wOuLLp8/yXGWyA+LHPDR0bdz8a1G4ZdKpsq
28VOeoqwPRLYnmKLylhNwihaqHncNldm9KMk/MQBohN8b5hb/Tzoxywf0FDZzx6LIEQRvcFGZy5T
v5ZX7pV7q3XzD2BtM/OIKytC7haN+PQLLyON3FhkKpuYpVzVaLKsuuQ8CuJs6M8cWl6Oq3KcsJK1
Pq3a3cHdJ6u1bZNYXKCVJxU+JUAJfWCcjJxDxt1+70Pa9OMAV5WhXJUT3yfn4wUOFPuBoyu1SnNd
/TfQOIeCB9ASGA/HEw+QusUX+JHdzRONNADr+cFP7wBZzXIk6ykICuCLGi9KFjgmEZy519ex3DLI
/qJW1LMiZl9nAxDZQZZbupl0LctkxztmD0u1ulLEQl5wW5RlsWtmZmJwRwo2rR0UxxYOCzoL0ay1
17Zyie1QAbzsNPkfTjc7JzAdMXfyd497PN2qVs0lhQsR82y6ssgUSFrEgflT3IbUFbMBg/Qdmlgl
K5RWc6NfiKv7e+Bv8I2JCngZWplmCFo+5n5dxuwyTjyMOh7G7C7Ru80D7uqEfQ/ZnFX9HUzuGsZ0
ykHP1XbkCqaFDrxro5Z4sABopJA0muP5RThRivWTsS+3grU0jOwXpLJp/7IfVAO0+MvvaGOUX483
HfSCovklyD/Gh08lrAwL4hjEY6AMQOotpHtdDDXwpoa7vl6h+Pl4tMA2MfVMUZyIqWUPELduBoOF
P6RDsEWiJNTMOB5UFbllWFacVgsfBNQkZq/Gfms8zm+khS9SUQTIQ64tFGvs0ixFcswzn76XW2SS
njgwe++AzPjwnZ3fy1fdlZlJ5Vpv166ITUL7fbLZjAeczF24NvxkrAmKD+mtNVNsAQoqCaya8yjd
zoDCikguqt4fbo/VDZdyodPvr5ET4Azz3/6kR6vrlEhF+i4TOXfWJvuz8uCPqSzqBjJKGjRFn+Io
OfrILXCbCdBDAwt07qUnRe0IhQMJ+17MQQM0eDu6k46wmloeMYY/erLoc9kAm4idNoBW+OnZKDGJ
qNkZQRdisoUdL62MckhoPVkGrYF6Ux8k3TpNfxHwIiix2gV0bYHR6XwpZvOSNpwkCMzLaOPzE/J1
Wgb1PV3LVx9sUSj44+bawrdvjz1mIgAKnopkHEKEsOOokHgMgJjMLdDaZNbaSzBh1j85emBFVAoI
h2L9G2mbgfHnzypo6K5W0n8dR/3A6lri+UTGdpG3RCokB78/5QbkCH5c0yWHb65X62Bl1cb9eqrY
YcGn5pvFVMJR7iVBNJrOOzlj+ABg8BTJzMrE1O0hfyhXLtoy9dc6ujBBl4KoX2wYVCiB3ccmcjZo
cM2EzWpsc5iYV0eUBbe/E9U1Flx4k2xSpkHU9Eyj6UfPGnFSNMYogZixyGv/hw3wedZPjCb5kqEK
R9h/IXkhCzohlOm2T8kVhxow+rUSzfHnjwl0pc97Ah3W4c8AjSmwcNods+8E6XAPaBd2Zz1c3hy7
wcTYhHD9J0ZIMcmTKFdtbi8LKrud/bTYbMnzqoL+bDnh6OI999yPyXUkjIKBr2ylkGsHCr/8EUj9
MzBgAcBPrF4gcW8mR/tKwH6nRXNFkAgBWZFfe3kPTLuK5m83W8rEhU9YmIJaczVfAi74mfNRyxGz
ZqCbfSNEdQvLMVtLKqEc4I1GstQtbtsXp5OWA6zLw+Rq4RhWfDJt0urI5jLtK72FZCmcvr+ecsaN
Zclo4yVZM7ICvcKRDScw//Pe0A4mqv9enhLyyZHpDnClCz+5QzjJuJk5GlIqogMeu5S4Vr5hziZ3
6yXrzO4keYEbtncKBm6g2RQfhS58h5EqobEPe6jN0MjKXob3QXo6Gl+rKSKLNH/WjkaPyrSsJRyL
Q4gQ4fpE93XDnbRBBX7UQCZpPDYtnjxhSLApaY6qWRDsCpnmpihNp6UMNkcMc9tMxttKw38Vld/P
kkdzEtATRHthHTH/9f9CAuGol0c8QUg34o2Ovo0+Q46MDerAuNH/WWMT7fMhOAJjrTbi09xBEAdb
PmkMdweXPo5Ggj9gL0rciJGAh4BiGLrjW1gWGCJ4aLbEkqZW9s/Y1JGz6q4+QjkwyHyirySHKDzG
dBhOqv7InuKvlkX1TzCJc6wrHnhETX+eVXAjyNvr5WPdzR3NcTRuTUfwcrNteuCFppQ9/ygxvblw
wgAQkB65FdkoyAwvEJgGZLBLMh14wSHjJIv2IkV6zWrTSjkCVdQ6a5IR9JS1snHh3y4cfzDwNIWL
E9gxG6RbCrdUBbaasbiMJDRoQkLDXh1iKoXKigJfcXlzrCKfPyBWON3DsopJAu7pLMc0vw/Ox5DJ
vIytye19h7rvsB0QPpMXorHguqz8ehNrMyUA/w+VcjAM/wl39WIcZSa/TpXFJIBb1cCD3xX3+zS+
nW4WFOL4xaTHjaHhHQ7a5C6kWCZ3+ORbjlZIb9rm/0hC52S+pU+nrNMr8TQgOwV9LAUdr1TsfLMz
F8mi7WRJ25/ZuKXv7K020DBpzN53jarwnzlprC85RiiOALBcOkav3RTBHa4nqRMXrr8oNhtgjYhM
8u2Df5KPmkVXxqJJC4nFfKDjLKX+7Gg8rX2H+WQeYtDxzuH8rR1DmvKgyPoB4uh+C4qRF79aPWrV
iowvSOyRIZN0ESohyjDuLJ88HqJONmnh5ukVgd8J1V5M3W3ZocnMNXoZe6uHZxAa6HSdaVTtQuye
wUzKW1UeVDaC4eUkhMHwg+KRVZQBOQgKu5LTBkzAL7W0qvZlwkoMnGUYb4QhY5GxRd1ez5YBK1LY
fVIpNqztb7pKniw2d5pYYgRD0GMVdEg7slhMqwjjd+GpXIJ07gE1leP+cULssGmJWRHBPM9DJ3FT
i5bjqzXzLQ6dzl/rxpnzIgE1cbJZVpDaPgqURMmGasEKp/2u5wOVgfYmFNnaspnxI4GZfVwvHksh
eRbicxlf9RIqRbg+09u5WEpoxI5wMvp2pI4Rf0Wzot2ceB9z5CIIkkkOFIHluBhb+Sy8EKtCuPIM
4qpdig+WIBguwzTKXL2C2FGHl24qQ3tqbfAXZVvk6tETYDr+QyiJSKEMAItvrs3qLeOc4wiJy93G
7r5xeK8ENe5/5iynE9BswSFeQjP/kzw23BQGYfIpG0Pwj8/nfvkLZReRT6yDEo4LH9FQwJTEWB85
LF6sL6PTcfbK0ajlLO1NzntOMOa6sHldFo2nHyn3IrIWSB6i5n6sEKNeDe/7uqFZLFwVCpMpveg1
nvx248fwzGiNL60I+W9IoR5EmC5l1Kp9IkhBYvAjU2rC7NSxMoVyIrlX+AjuI1w4vXFOczA61nDf
DbAzxlRDFYbouAUAzfqdnKWeNK509O9hlqBezJTPn370SmkDq3Y3La6vgKUfsLFpt60KjEC1k5PW
XBs4EmLuoNl7+s6HAlb+sBXaJA2y5v+gi4BT09+MbgBZ+a6WNGxr9uQWO68XQIdqrTE42Fc03JZJ
FQjIuVpN0n4ypjWoOhgeyt2yyi9QVGC6FM+rUFmJZmVOnLs8ppWPZYXdF7lh7wSCF2ulm9Zt0inv
Ezizem/qGDvWwaYU/x7GFmxP+Q941f1R5hgau/44xWwZVnl0CVdloGQCbX71D/cPFaWKKYjJK1Dn
Rpqy0YJS8zZIh8wfBklvAIbEroxCrc7sLt2s9squk0BqTcjmUUpxbuCu7qJ74D1/WpqnDLzM49OF
vJ6tTLOb80RT32MimbyFTXcQyJ4Y6ceGZrXoUHV+c2LbMIvfD8Cmx2tkAxfa1dazityZqTeOJh49
peSLyGh/NCN5fBCPD8kMlisb9ZdQfdXLpmv31CgAUNojeXylDbDmAAhwHOugvgniPYT3v6gddvnt
flICxcMva1BxScADhLFjxhNBn93/bUGCkFXfYPNIP0j4N1pjtkY8kirq4B0c3PjxtF35s+P/kf4q
QWlbEPZI6/uXqSQiDbuc+uBNEKhg2UlOzS7UJ/cQuvGg7NBMnlKb6gFT7PJTM7Ixb0o2u1q86737
djnmTDsmCBrgMgz2zwA8u+/U35nsLK2BTUxxCtEOfLSsHESt2X1iACotvaYk1B9D6U3AoStHczjq
PU9/3MVU/AbhErnDDQLdJn7vAChmQBQAVJ1g2y0BhkJ7yzAp4bfM/NW6GivEo5AllzxmSt4ea1F/
jWEw225HXWCmhm4RiGkE+k8vMXLH7b3loc02/2cx0zTn+ydJwVMUNvS6JMVNgviu6A8FRdAsVo+8
xXmNcK2df2nNUljoffrfKXkk1J/NCOu3Klr57PRD6y+iDv+A79f+KqC2Uo8ZQ9vxABrZWRMZjWg7
qZ8b0NUMDses9LScqwATIsikC11EAQ8IZUTURe0PCE5iL7KqnBtYLe5+VkYZkIrZJSKESzTHg99X
NPLIOb3nLnRYNIwI0cWoIV/sODrgqEZ104aiCFhnRkfrYhU59JG6zv2WFzJvdGXa6HsZCX1OtAIT
ymo2kLLssZti4vtc8Z+W2Dh3TXhWhmXEbHY2+BBTZHH+zz943xMddFmsFAZC2ob7L7VSeGoV3C4K
9ZnlgcuXYj4tecx6zHJ61Fa1oV7G7LXwluRvblvn7AVoenNXPJ6Ef39gNEaModl7+qOQs6KvNM1B
LMdLWG1a4cZxmFVDszoadjpaSPw+psfs7+Jaab+HhCnWFAjzJxIRmldUTfwY27zg9N4wn7FyKFaZ
kGRyc326S2niV1VccyG0nZ9xhJyfC5T1HeNUrgQhl7dom3GeIRESRoPqye5SZ3reAcKXJA8Stqj2
ddegSQDSx7bV4yYBMXZRa481ak5al4qZ8EhbpSx3JXWoKXgDpfhFgYBY4VU/gDN79jIatG8sHG5u
64oIXQaLoX27DwmU0HeAtFgcUi1tW0rSLpv9o8uSApmZhmy1QC6Sm+k6mhjcEoeCYR7HgsLHyQS6
rQq5oau1Sty65XXjDKglUJwyt0ZV959OfxHJ7NRudUxWONX1Si+/FQ8+kC6L9TOzzqBKX/v3st3p
K5Ii3JafUrSB6LHl9q9RyTPc0g9lKtGfGFnMw74uGNWsLRn99eFVX+fGesl8wX9DY3wfy+JdiBfM
Usu3cWxqii2fch0X9FXVYAnKqlv6KJVsp2v5RAW4JWzHwoimvmBHErDNHl0R3SdYVcJKwILmGJn/
Fy4VAdX8lnwSoVHRsVo3kjzrSqaYsWIeyHg2OvlWznjLYh0KP69OWxNrRGIFPiJDD7r6FmFLfCgP
mgF4pfyBQ/0uIjlMIcMT1P1wB3UmGM5mMldL7BMod6e5obF1kiC7+I557OzheZd7jDFf4XkXcRH9
7OF9hRJAnvliNyKaAElwvrgMOFJ7wzcOTwWAZs4lBnPObYrGG2MkgH3dgYtTxAT8g8jNtz3ZNHV0
0u+R7LLY7/5rkDzoYkRppgOfFHowaaURXVzi8NQj2R1JcPlQ3OOqySPiLewtl0S18TjwAt1YNst9
5HApiSzWZVlarMhWpXSeP7UgrQKY0TGVf5PZjINiHqFV4uwV3yenMdoDjaiTaGgas8hZqhKkfP2s
SaHPaXNPeswQEYzx2XIpxaql/FVa+L8zdUN48yf6dvz3ntqHtF7FeU5PLLVMJSBS5XCW1Gp9B/mj
sxONfbp5lPf+JdrPehPIJSWJXs7iZ7mX1hnWXIypApEEg7TePzdFfxRQPT0eykonhUGHGZUl/oQt
Zwd1PtKGZ5au7fnBFOLuZjUibXunumTbOaK6/Xp5ZX8vbYHZaptE1y8aJr0N4TyPE07SIse0GyTY
7gLAv5TgUjdJSM90pD5cOGHTvTU3ekImAA0d3RLN12nJv2KbTLTSfcP/5+uiwiVaZdAViEHalWIf
rtS1/MiXTgmHuvClBhgQWcw+KTR75a1N2F8pvG0qjMqnRQGVlgKmTNt9qLGEjYyR6aOJkGbkbe3m
nZRMRDH2qLi52lnLh06KXxIoz/YPK8Y1qegInYGYk1aSzsjeqXRnTiS2FZ3E5AzDefRBpulb53Xi
xyzXHrQ/j1ozy7M4+PDxyyQVedJijXeKM2227mtS5tmPST0ikFvN1ltl+EOEX2yTeouMMxc3ZqXJ
Mz6W7xVG/mo9TZmPVJ0fAjrKTDR2i+lPM04TFAWpKj89ONyK+chqdwxZC4TdVYNOWrVag9acocuP
kcmrtEolIssdA9+Fp8jZ96aqZ6EpVMYFNZNVuW0ww1Dbao474QzEqCHuDIBbCpqUInlLhhRr90YR
psAqjUDUmHUaqH2WF2P3nbyR5btmzKldzNTULs5zpxCbVZH4iRuGd46ofN9ssHo7sPIJMuNFciyC
QpPsvBmGcPyOo90EWt7axLzBOjeUF4CdfoTJ9jesxIbl5XDOBCUjOy6DacnK/KKcDgZlGCcLzHoH
oew5gvC33XdLo+E52koGYMSuLgrqd7NCPsXewnLlN3ea5Ea/dCj8CasvvHYxM5emzCqsINoMs4e4
LF3BrWF0tg4Kvd7amllv9/upSeytAQ9j+XWnoL+gLQq8WZcgPrQnpK++D5hyS3MGbwEZJJT2MfMu
Ydpx7n7tO2+AAqtOvUSAwQ94JiSgHTVA78//MF+JhSEGTwosO7WG5y5C2Y/O47Y42/RMqVsu62hE
a8uk/vdCOl8WdHnZ6O57lY7Z1E8Yam9e1miSQ6WdSCcsT7uWynRb3sAeAo3p2fJwk6bFjzwPTtnf
Y7tNtTCQFBMaAFvzv7GK3JdgwqSOGc4ulkjZ/F1EQ/TGAFJv29yJ7mnrjD9HM6/P+XnO4hmZg5+m
jT8QJIdSuD/RNrgaSKSDSAYnq3diGj16/3UIVPMybm94ejGyPlGn4vH4P5ajnRBjdK8/1zA/j+B+
0F1/rD0nr7tiMIcd41jXeFoVwbMvxyQyoaN7LvrzV5TyW7z1L0oE1ohcYuQELHxiGIgVSoFypugo
KW58Tz9cSmfqGi6LEWPLRYq8667TjKEGO+H5nZ2maKXlfVFAl5fOdN/9qmTrqz1sEccs2sgTynAv
8oba9Y4pUUeQK86ddjVIvJIBeDzdLsp0fY9DQDEpOj6nHyas8NxZNu4VY7Xw0C+eaGBJ2NVbKNjl
VRm5L+49lT4SEsFzmsUAeM6uw2756fN7nG7OlPwjeRTfhr9JJ/6G//rfk38q+o2uFmn20mzeRsnb
LQNODvEDEcK0o09087sFWU+p/1zLvJfDEVbWk/0hUFKbnynwAkhl8WwiP30LiPySyM7qj77G1vYo
iSwMUyGDuMkd4W0AjZCznL/8ry81bt87tSEIw6M8Oiix5v+eURegwz2PgTDh4YW6pxcY3wCVXFEW
tgDYTQZY+tKj2UDZvvFLlnk5UlF4nSQThNB0vey951C9NKZIUZOtxVjs5S8O49XE8EdxHcszmgpN
wDcWEUoZvuo+y1V/tMYuJKsEzk5AIXkr13lsSdD2GtLrG3j0B358pn3ZV1gyNH/48NbEY2Yr5F96
S83x0Pd+lcMm9PtB9TU+wCZoCZrEVjVo2Dl1v6MKH348p/eZekwyKWA6F/G66kn0OhPqGxbsynWG
9NJZhXUfF3XOJy2aiyJhpBHcFbw9TL1IgiNhxFGxo49F/AlPGo5u2ZbNxBtX2097by4AEPMzGkx1
7MeWnbT+aN1QHPLZtfdkdmb1tjvIXCT0otxzNcm7d2LemOp+2kbylkomkdbzCYt0dIglqTaXlYEm
QRCwEcfkD31mKSxGANG+QqqSkE5C1BNfEHJEIdDfvB3saLPYhtbWFrbiQlTnLjb2zbd7d50fmu0H
Ig4+VwlXbRfjhO7+pcCTN+8YeKVfUIO5vR0ZpVukGBC0t75m2zUpBhlua6JXbUsuMiW3YcjbCWVy
v8vzD/H/T2T7c1v+9VdHJh67SFXk90EI4JDp+2y71bagSmgqs/wGB66SwLnrqWrreHhpS7Mehnjs
7CLA4n7+RKeAvVrtnoKxTiolmin9CIjI/fuq2WVntNFcysjTBuOIgJnf4ZRbAD/yjYY/W8oURVBd
W2rB2QNyEkmLepvZRnkFlZx1zoFsDzMYtlB58banpLMfBhh4jTyZC5kRGlLXF4mQj4dAE1Jyv/hc
1O5bDWg5yJzmS3igPTXFDBaphUvpbFgoIGDsH3m1nrzr2psy9y8iK4/AMio4BrTLWSV34jTOThcb
yeP8EPZRkq2SSsBD7haFw3y+Z6yue0R9ELAdLiwDcyh3FGFDmfcvHrwnncCaQBP/iG2B4ofgXero
gOe8ysdEtZBYVPxxBMTY8Grcz+yV+p3oyPmCrcdVRnHMoyx+q8Muj/OLN4i3LbULGAV4PnkfO/fI
ffUfXGVFO+YQjDQcxJWN7riV+oForb+om9A+WFdpVM/rJ8lApkIndnj8mqteP1j9QpM0k3XVzloy
iR0s1vvMp2bCYvpgl8gP51jLS52Sd0ZYBnsUdBwoE3eTvIgMgaQ7//fAoO9zq4JkVp9m7xAKsNHv
iSYq/WHs9VUkabcX07QhJejRn6NTOZX4VDNeW99pL4NxOIgeEOJJ2L3RGCZFGT3y6EftZJqf5EkI
HBwmN6DTnkpiOUjAcnaDV7trdFKpV0PH+lJO7ZOj5ECGBwmzu3JX6Ayx3cNKdQsFGG9Qs6cC7jkK
2DBE+flwZpvxW8h5+eT1RWIGtkPwOlzC2VVAx929ffpX6Zk7idjqCqJWkSL7STZse6Vq1ZADwBXz
X6ZeZWPavbsjT4cdukLlKMahmJ6+hGJvCxXLOfuL2IVcMyH4Y475mPH0nKeZvPf5HImJD2WNgIvW
OG3VRL3Hxx6uLAg3UFZZoob26g8WnkucYMLDstWApuSwbLZSXb6P+4PmNJBSD5YmLmL7OblCkMBY
dYyV3953HgxudEpkolTopqXwkjQFtfNnsFJowcMzzevYtsL48oUE2Q2chVWAwMAYBFGBKoVLooLR
r0I2Rxe0O8k+I/FVd82LuqT6IFWcuhfZxb9s1aCUaQBj2ukZu8NJuhNR34p1OSN+iQ0pnD9hqUhy
LMH1mZ2G8i4zZbvPw9I3scfvNm0xTQI5P09f03gCjRdMJJISAnx3vMG1mkNd9ihFAphEhslJZ+hc
preZQ8wzamECDdiTddrd9gNbBaceS/96cZPNLLIctajVlBctQjhgdy8O5bmEr6SfNtTx5XUWOEuG
fWDWZz48uBPbmgv5KMPYvXOdHESD/mmflV2pOnAPInJuw7DQiQ4slyhXOKXsCv7qektYpvAt3nMu
7kxKWGrx2kpWo8MLo0T9lDvZBgkUp0+YkR4u2n2yaGS/aoxRJUihX3dCd9skPW/zDZ7DHLi2q5s3
P4oGQv4Xeln8Z8QIa6pp9vlJRsUrby7fl9it/+CYo6PE2g9+FE/1a2u4isnBK435SZg7hLGJ90ca
90qyaHUQoPvdSLnoSL5xdng+9ugfTTrv3XF0F9KhIGEzbOyBJ1TuAxJtXz0qGnH0oODQ1D43CUCV
PwH0A1PDMpdiXcNV6yNegCgy55qgkwSixCOoQVX529Ma/2fiwmk1I8YiSFR3baJXT+st2AR/BZ5r
sXlT9kPdZx2906rBAkEJDIbXBkAHx3P2dDlTRLllrI47scmlFNqZGAPcZObGhJsndjsyYdXVMTR3
dkKYEq9/6FK088QKQpNyiR2KBubHnyouNrxkxwodiIKsD9eg3P3+J1Ob8v1sAqNehnnBSL5D1sDg
kMqIyby7qzD/pvf8v4QV4vmtidghR17OI+FmmIOTDS+iuOs1fIDUXJPcu/D5IEsIxG9Uox/MqIZ4
7y80snyqUG9MU46PpifM+SiEXuMn5iM0gM8cLiwOJYTaJtB6EXZLu4+U3AVKypGIgOOMEFmeM1q5
eD0PBKnKoutrVdPj1pRCRNiJmIb9p9MSFddDzWlv0YlFk0V9m+G7da6VBT0FRJYSHCiNKxq5dpNo
pk9BhgCAS5lh+VIs6GplSvXfJ/QdAUI8s0Js1csfwgqaBdeO/2rpchmCIHWfWdamdIrPqf5O09tQ
7QRdwfPSZO2LjeR5egPwjhrV+UGY9KJhu4PZsK5kkhm+snjTw4p+sNT304anAHw3nWWrKg7QPChv
wYtGrFbuZjIWLYtBk5DZ+dAc7un2Qk7fxoqJ265voBFOQVFZxyxFXSIs/tAxYAmnFtmUCivIMDWd
8LExnnuUxsYz7nYYskvhErHR4GBsmVi9ShnDZTEj4ilcIoRmgK8Ln1ilwIiMRZPknijh08plrpZt
KP1a2D4WCk2TQAsJCL3+3EIjUVplg0TqC5Ks/VjpSw6yE9ryT32FtdNoAe/vj2Fw2T2x1NUuryyv
WkEmJd5nlCmzDR5f+nwTORzIkiravhjy1+roEEvmD6/SewENYLahet3W16zGeoGR3+ZM19IYShrI
cYFz0BkPdXFeN5MERXQ+iQHmJmbZYU2HokXG0xVfdNY/FxXFFk8pOBkY5a1DwXbA4cJAspqyRB0c
PQPiY3Nw1qKmz28Ndwwg1UD4/jCdOEh/MC6RnwWev3gpHBZcYj4SYbnvXhPpOabe2eqA+G3qCabP
rHuSa2m8zwln3EowHyaJ0O02XeFaG0oPeGdEAYkhqZw3ccJcHBB7DAwz/ixgKLn08dwkRmbIgh49
rmlNOm1X3rW75iUIQ5bmDdwyYijPM5uXqdeBl4SZWnpEvhQSi+mqltlC55yDOFL/XYEMzEG7vLQe
YWIGUp4mPvDvMdLtpS+1IiwXWuRRp0lSKsQtoxJvROf3MRibQuf6tyRmKOyH89KQEWdSg1OFMpMh
uG5A8jR+o5rZXUfaaOkgMqHXmMaycBzr845XBUGvb1nfK4jtVe+UG1N8wl6ATEtRqLrATZTtEvvU
J/fQloT526Tdio3x9vEhgLmMMxrSGqSS7H1074nTzpSwpjxFoTdBGfEmO3eO1IbTjVOCxk+85DND
+t9rmcOCycjP+9uZ677CIcYAgVT7rmHN8Yy7TtyXcB6IJM1nbXwnbk5Hmz0WP1ORMweKF2pwnQRz
XuiyTXELrSx3sjgvj2H616A9asgzEuq7rNPNwRQl6aSI5hexwASeGLg5ULQ+4h6L58bwU8VHGa5L
5yM3e7l3CZ/UqmRT4WRaQtC9epMyXPr5nvxSZyFAsz2Wgc4Uoc/+1JMGxTsR0YrtIxC1u7M1cQbx
deHtW3+VcZo3zmya2axiEme2+HD/na1ZDTyzAoUyOYoTXQgzwToZzjP8ybdFcvekQhiafjRQoXIT
5A1k85U4zyVN6ZwqRPiQatFSJJDbpFgjlv+oe3QMapQ+oH2HKohn9ZFKlQDHmX+aVsQeEcVAp3Xb
czpwgI52COuYLImuSPwGlt2S/LLKA4hxlE7iE5C/DJmfF1OpXWo+pjcu/0fqRqUICUFGlE9t642Q
BXDfvAF+47nNlfvYF060HIs4JC7XZoGBcbhLhFGxpuXoQZ37b0dRQE3/sZS4L2hQ3uhRe6/INUb8
o+PHzIo/uir+l6zzjWI58E2Ao+A5xS1APurVS7yhUgPzxzO33sQVpazZdlFMW4n4LvCMcITCOO+z
t7Gqv5j6ycTOvsxGXDzJYsuOkP9vK97ozHxi0m0Cq//r+SqtYKLN+ZIXNVZyVRSwuhI8qvCkMHVl
cPOyQfuDM2KOonHg+YXkS5qwxiCuW49oW/SjZ5ap5QRzBEYH6NkoxmMYLkSfqv5LuJy95K+u6rJC
4mjrT1+bMsqq4ekqM9n6hXqZ9nB8lq2YKEZFcJZPlQjTCcmBUK7KIdzgNJQXi5p+QgrP82ZNTOJb
m/W7eEGtPIAYcGKyR6ia9jlOtqgfYpUKjBQ+q81vrP1Z/V19/XZZvSInBoPr2hrf+9SqtdaZsWT0
2SlES8Jz/5j8F/Bml+aff7HY+Mk8y5ipSJ549ARSkhw5tDJ092uwrUeopi5q9Fr8nvQvblff7SQ+
hdyj4osfp0JNdDxj0KOiGceOItNe5tA4IhxdWx2m7cpVOCZHoEi+dRb1exQ/ZB2WsEs0mNeuOzDe
CA5dfGASX7QqSu8CdjomXTQ7AozBSfj/pDGtTlD4JjqvL6qYmDQIDn+cNRX7HFd/62TBylUDnMcF
eKCNmh8iBpRwZo0pepG/ZIcU7gn1gL5pKsXv7f4kM4kTlaSlK006HffaR7yZzilc82/ogaDKjVKR
e1kt2k1wRh1pAT9sc34Y0esnI1uBEd/7QWJJQnHn9e1U47qGb5f7l1cl9815eqVZTl4iYOPrH/Vq
6mY/Je8Pu7e69CLvJLF18FXyYqn0+0mRVnyMvovYrAkyLvpZ+k7D3ssfc/TmgZFAAaj9So6s6zil
yqyfNoMIto7ONWJ3NU7uPxOEd3HyMIpM/WgmTGL+uHQSMi8n+zGxA+ytEY0t1dDERb/kZt+Cifx3
+kjPkOC/l7LPQuj2uiQGn5116IZsZ5jDhQ+4z8w2estq/BEZvWPwq54+ztQdun1tX4E2DTcS0BnN
UL5Ew7ZLuwh+9MXqHAu1b765HBRuyY0DTzfvIavC9w/9jmPQ5rQ2eYwDILMLudCJ5PGYXX8wOYWZ
vpyobp4YqTr5RT30qLwUqvSGIbYMmRd7SQWW0V2rJSCz5P830ZN3yl3eXSGtdC1uWyLYs56POspV
7hsYzlxlJwogC90fb7bKanQ0+r4DdLZ0mYCW112m+JZ7U1YxG7kc8Wg8JZTmXavYtcQwe6ZASs69
Pe2kUIRLv4WYxrePcHMEE6aTo9E1xDoLJZdhKIIK2Jz2and+6qdELTkAbuCyoRA6sveXFDJRNIBi
ovs0Dim1rrV4gczm74+EoOp5gy5kgg/KaFct55JOIlSbd7Lj6aP7QHgrZNVgmyadMZ64PTZOmviF
Pg2zx0UVdhyAigVsCMLspW1QApvWxFRxEFZaaFaa5g3GGS3Kmb/Mbqr2eAfz9NAU6IqdINZzSf8T
XLThY7Sh0mbg87XTezEqI4CvXcUyumaveTy+lgOBMZCFIGn23Kt0kgxZDqHx16CiEILi8tT/kWX3
va7mkNvOetCKh2nzH9zpxFxW28/biNlc/F7TtagpZ4HPsvzLyoKIMFA7PsTa7zHi1O2xvdthUVNk
0oZBSq+P7sW51vV69It9SNciwz1PKWBBwl4io9EP1hMkStAKP5nblSuJq5JE3ACovuvcemM0k1j2
7NitxRnWaqb+K6DpkWDCOPCShHZhfs7N7MwM/e5lJA5FaQjlELnqQKmekPQeP2oPtbnQMbaNaydo
/jlUgd94KZlJ8NHeVb7Wx9sYqlzhwW4aaG09fdqMVN6+OONuDeeHSzLZ8xWJYXzDTlAvgxIjd37T
TY4Ky90RiXmi0oa/hxJR/yyNQ0KAcOWnNnGSQLTgwlbYiRvb76cYeirn8zH5T1HLjFdXnhhvMp+2
pyC7+bMsfs2CAsjNbOqF97fAdbHcnc2uMjdByYe51iWs2KhNy/pK+FnAfJVJ8ujbmDaMMqmmIFR+
9VwtcAnMhYJXFcjauq8hS5d8GkF0Hu8RvaDsIgEBHn2y4xBMM2iICFQRAJn3OBPrdjrgo1EOLihb
OMLCgpqEE9IPyXO6avPpF0R7aDlwK9T+XMV+SYj22eUSfH+ZEP7prcxLsJK0yBmJ/pLJc2+BN0Jb
VZEePRZS27EAGW6T7fcKhXXKGdt4snBz1GaCWxnRypvbGLXeiiUNbZKcu6BRoBBjRWnWFMK12qHp
zZIGcteeiiF/KMSgImkgnYeL8OHgjrMe/aJ0RDY2GTZgkElF8W3c410bePJXlAxAPPuWG34QjBpf
GFxQc0b/nC7QTdUkkTw4H6z/wZUnYZC/DgBT3fBoQT7rVebJx2uNQAdg3wLa4QfMiwOeiQ/saOtY
hztbw4e40vtf+8XEOOupGpEY7jRZAPxHwYJnocEaLBmBT/bMzLIZtb1Mvb4tJeBiLYFtMY4QMMNj
xMLdDO/d5tr9mEkxqeiIn4DPb3xzS2eEr5+1/fJGGc1rMTbHV66g7ePpJUag16gvg6XJX2sxrdAE
qFiTSlaxIZ3Siqx2wXchKuPsNUE9brki7VsNmQMTuxqZzMvLs8JL8BgN5yp700YFGkD/k7VX+GCm
nBu0T5Bjzx7ztRhhlQ5f/Jlr1chLKajAb/oThLyxRQ5ojvNc7Ds530XG1hVDuOrQBVFIZSefyqSm
51Na40mf7DiAK0/LNoWVvJuyYV5IH4aa+0wzADkORBDWEDvR2ENvQXqsD6KDQBlTFxGQKzRErt9+
CP/gjotTA2zzf2eBnW5PiPRf/21bQaM1lgGsgQMlvh6R7v9sH+USJQ4i1SJLx4TeMqGMa8KlKnDF
qBv+hfSIkVYGEH1GT6d59D1KZRX9eIJ6hCPuWXQRhHN/HBSIuUDixidqksf256J6OeEa2QkBa/ug
KIsMWunirQ4ynxHt/MRGBXpTCUFITSiThvBRcTyU+F5yZdJPbjhIrLQ/hnl+tCo2vlKFBJKJcE/B
WIAH25vvVJoVQ7/ydQ8X0D1bPR1CHpIfmysZj+p+9wB+ccsVPPkM4iPAEwRAfVrr/vkQpsj+GTx/
4eF0ek7s5wE2CMddAGTE8hQhinb3yTVKH07XHLSuTf3CNT3Hw8Z28YzTrFs1RwuI9tn0FKK97q+L
2Om4P9hV62qWgalrX0OLBalEsx4mq/cKg7HbyYHX6cfbh3sBvYeisOTqJvVXQW4AeFtrilmwjzJG
KQUSilLK1SwqHnifucOpVCVlcWx7yIvIWEv4JtKHZcTAAS1LSd6LnKbKwWEetHYSczRHs/nQfRjB
7xNxe3E3hANY/4tQfaDVMwn8K/4P+Gpx6IRA/lmdcjZg0vzaCeVmE08W9IBWyOpntPWKv8OLljBB
rH9SPGrMpiNIZyW5S2KdFZhODdL+GovDet22zWKEDUOlGCYAGyd1BqeqL3C196Mx/8leEVJBl+Og
7coQbxJ4CZjY31dS+cOBFzgMY/DoGA/6rGfKHAtL9UK7iH6nwDsSV8KbWn5jkyefFoSsO/LdhQqH
KxqpAF2op8pETmCdYBUzKNpMTx+s0E3Q+xJnzFOPqvirj1dQI7fF3SpJ8WipeReDK794iXa/kjld
BBGUOusgCB3snvdKMvfoYUR53VtANW5oQg+PO4s7/uS2DBG0JZPjXgLe8VzoNvOA3QwRQxJC3ZpK
uY4VxQr3wf0z4s8p+PeDLdV3GpKC5DWLvFGiGdGtkz6Orp8NTKFLiAVLlRheGxQdyy0fNeJXePrZ
ktbr5AFhkaeJesROiluJptAOmxdHRISaSppAVOM2Iduu1TuB02mU3UUImuaXsjFnrvY7SBQAnUxd
oGWHQq3jJGLqpL1K/8KlZK5D8rT3jcOfXFiMmkgoTwpxa+RuMIkdi7JX6vP0mKAehOE5lhzlZzcx
h9lVUp1qXQz/FNDYG3vq4ehX1EJV4qrRJcCrPOYPxyljT0yZ8vswUuj5L5ZbpSVDTXWKxEdtQ7pC
lcTPOi1+iYas7s0J5RhYiRPiSp9AWDJVVg8gpeVeShY1hrNvI6UJ7FVL6fm3mmuH3UA/qJY02mYx
q/rDlun0Sd7A6NSLMfX5n59f18yTCg1MIe4OFOIFNrKAGH9c7JuHVPqGfBtCz69Bf8NMBxXfExUS
L+apv7OUoyKDR4L/p2S7wgq5nUdKsswufD5UZgyz5sObXoZ7rbz5F6oSQ3xUQ6DqPNAOba+4Zx2y
NvfYRtoTBK6d6K8nkc7pQG70PU9ATKe9yME7k6cfOV5EkENM3KIy2PZKhyki2014+2bAdADnq1rx
DukO9tB7IRByH32m4jt8kTcpK/CNxjhwx6tJ4Zn3KDhfBLvitPpOfe6nIm07D9PqwjKgcDAWmmpY
hZLIiwv06YevqSE90BB6CMzcXEBQjSw5yg/khNTiypWWsJRV9IB+UtpW0NFEkCVPQAaWf15q5yeE
6TXopo7D7m8Cam0BrW21Ltb4lWix/z4h3wmULyjQDU0oMiqHl6TPHxfNPgw6NPwuDE++sCdKyCPS
z+GZUwjLcVyeeojn15nBV6zlAvxTjeQkVTE+/f5XUWXMvM6KgEgGOsI04ldmCS6A+0KCi43x70ki
4440kVCJueFrny59bL2SnGDv6O2K/4+NXlsqBCgBT9Jg4HbS/AkWRRHQDCeVeNa8URYm/Ax8sCA8
t3nO8OFpHgST4WcZgjn5DODTQOhv28NpKoEvjYoGfuP+c8E9QnqPHlVzLfBHZ5hYFhR20h/5xo+A
+qJIYRGZkkCqVrjeXzKBmY5Swaa5qWM8IDNWPs/mYZqQ6UJyCg+pUuFvEnAyNleigakDLnjy5P9S
RVzX4mjSoo+niPtOB7oGZqGZfluX0YPFvKGPjkPtzG1NVklmz9SLwnNxouA9JVbTfTxU+kofGvSY
sag9aNdgYBouxdnviG6HovuTcobdoCWqL/R5XGLXZVveOgjOhIUAaNe7WmwSJH8Wj9/lp2GVqO44
uICcBlW3mfON/Ox/TtCRs4y77NQ/z2wfnii+nropAvrhffCMW00m/QkvEam9VmX6HhhYqSrNTz82
oiyskCormXF4DqrXHuOBrwNLGDNTRxcpgnGefkFnxeQkJrZ4OJv7x4Y/HZ9Vv6dpacIGFoXjbuA+
K4Is+alHG8GKLWFuPNrHblY2eirvTfRrkdAKl8nlrbYLwtR70taK6dxXDPOA77dxRtBqZhpsjpsw
tG+JFB+RzW+RfoEFf03eE6lVNzNWOHWidizxhytrIx/WBNTiVgBG4O4VllP+gov/aRw+yauj03uJ
DYwP6wsfPcrZ+qoZ+JanRWa+FFPfICk2w1RvLugPXfIun70wo/3X76XWcwAzfqv1zG13s8vLkRIx
TeRikquz/2SUiYyVUbMDqGXRuGevvo0GGsIWuKB80MWQalUKakcPuQVwcr+yCea6CYynkphDbGXR
i/ewrftkiThtwMlwYr8ouXlJj242e1FqpSC67UKAhdLlWz/bAbD3jWXz3d3Z969UOJHZ9zwdU3nX
P6otXepJbFjIFJy8bs3C2+ppGAKTmHf64MK0/UdSBPPXawC1efhrd6ps9gsgIGsrn0onnpSZIBR4
MmwHdadbxnUqxrYVNlWwR8jGKTR6Jccl9J+bpFABWq99AucFBohIts4xVGsz+CojhV7T8CkheTX/
azM3qLT/bTlL/CTN6SPiwaivlVx7ziTalEN2nvMhWa73WkI4ZkfnElkhL8Ggi8AdKKpXPuZEPMRB
CzhLPa6sWT1BwU+DLHUAeQ3zkaJQMecLxkkkG+BbQtrVW7rvf6epZAU4nVVz6tdGF3+LA/hH1KDe
VmYUu6rIgaHmEllvk3tOGpvT31lgNARha8BrIdxC53LWV7ING4PKniarPA3fi99RDjHhJfE70bkV
ZqE1+U95JPXtFSQRraKfw7t0aHu5gZ1Hc1AuxW2r7bN0SOscEFff01suXBdc+IYWJllM4jUnhzbT
XpDKrE6v6dSIJJ3bWyrqJBErNQWStbnyGk/IqVYIifnS6lTV6KDcy6pbufaM2DXZ/VoFk0VULFYJ
s9JDWv7jBCknbmkSapwL17NhFhehxnS+iut6fRLLGG+/LW+FVwNG0rImBPg7rfiIz2ZTLDs5E+uR
p1wEI+LVxgzFNlXJDGKPTYswiAEdlONcBUbrfw73+rlBvk6/BczPTxtwS4J+4gpS3K97/EcDfMOb
1x7WkJzNjfn0CdfY6Af/cskYEzviVGI8Aff30lbIakapIVjsfDnYrMQ27JyJze+5bSldOI/lGrv8
/u2sNeAhMdTUJQp5Ew7+diuiTQBtG5G92uBo4WQmu6pu0La43oNshLsylQS6jUAVjMK68TXnn3YI
kj06jW8iCKrlbriD230KYRm8qC2CRjaelGW+HkcdmOVMXT3x6iH90w7fVCTJcmAL6n1KpAEaYgR5
2Eg+Un03EBLDjGGqOIcnwxcC06uKhQSHjr98QTjjQxQ5s+mW4K8uzCnNDMXFnNIP8E7GxrKZ5kLt
Ch1O1vU0OWV4cGyLm5Sn6vMMLXa9oqHAsbkhTXnKRSSSnlJIMzlUpa3YbHriUOrWv3MFESD8aZXd
UuZ+Jmnph2C8BrCQCcnFnphzwc8UfpoZwOU4XU2EGJUg0ZScRG/Dv4Sqm6whjOTYp3YbxkXxGt7y
mFpR9yGsvgg7YXBPjr2eyTeViJie5Ro/L1uUAvTyqgAnN+QgqkZv5nIQYEsrZl64N7wysFDCkUaC
pDNSukGGOlNsyFVxvH28uucX4jN6FSTJPmy0AXXp/fo3RqLs4TgfP8VpDzV+673TqHJpdfnKKUYB
KJG+I3GM8DP/22ezywcVVhKt7sRxVgyyWfX5j76UlbLDrRqxc/H+giFvytKaxgp1ipaFHLguhlu2
JCM8976OBWu7X5YRrg8jRI5gWi3sAkKWBIBgnHB4IJlt11zhlAF9T7YClgmviQ2opoSHAgVK76y7
wFTWd2hbcidqTAiH0w5LZiutJQBvTDrmQJvarfrjLyusQo1H6JnM4G3nhcwT9gwStQ39sJt1vvR+
T1bEq/WIO1iPklLTdvej4kVcOiZQfPuIdrYi08h9yeL/nkAKwVm1Xfd2+3BWaEB9SU9hmEs0Ehgn
rAFaSGjikdeqf0OrvdRx2Tx4rHaM+70N/pgI6CPC7trQxZWex68Goevoi3+svzrt0TfZqb+IZsBI
kmeEk5/8Ru/G13grp7AaItKh5C+Uik/BdmW/eNjdplPwfQW/BScUHj9bI9kYBTJfRr9SE2LOF2sC
ZLmWH4qQH+yabk7XkI9gRrS6iPR9jlDx7DJ1FzUhJ++FL3SUJjtZW7XrVVdypJWl/gNnvTUqxSh4
8W5WSGU+Z64wnzb3jbLismyrdZLBm8aJ82kIpqrlnDUxsyTuvZ9JwPv3f/VHVxhnR9zu3FfbqOBw
62UvBCLvjwxi4Ss7/3zzwpnMSDcRJCiJUpFOZ0ZnSj5sRQbPBQ+sVfFtnu7JwbRQAJ+nS7cPxGoc
8I22bq4VX2FgkaElknkgtqHh28DizT3W/8ZrjIIwC+HCNkJhZSxARP4Kg6Mlkenlo1SrvHJ9jo41
crUryyp9Qt3O0REptemF1mlj1r0bez3ltr0jZ1Ot1TDkcML/Hr1wY9Wy50gZKxDZDoO0Zh2dsfPQ
v2m1BwO8wAhgjxB0fZlroU5WqQ+QM7KKVJ8y9e1Im/l0pC1GMc1EfzNJcIMRjVBbc5UMMxf43CEr
Tfxix7XaTZ/6+DXXO0CPGDYBZguOj7G5857BvveECoSHZ/wAHHRO/tIJb8LuAP4gTKk5PNj1Artl
Z+0SntzYf0PxHKPqvA36DY2j337eS6HvCt18GHpArf+qQ3Bzfj4XibsxTUX7NXIavXO0ah+Uj7Vd
LUFyp4lgJDxzNxHrpg72EgOwa64aVZYn4vq6QrhyVXjfgrFkplbljDX3VFdYT1sbzPsB5IGE9qbq
SfVp8QSc2z74jO6eLdvxOLZhLM2pzt6D0ur+Rhr0xadWR/ZuLrgsgIqTcvzDvL4YUR/vasHgYA/B
WWn8kt5njvls2Xnt28zWzTecUiiFVc/Hhfw6/46xjN23Kc9i4ZmDoLwIQaXMTBrMnQ7I/Ws6OjZK
UUmr617RxyMlqtLbbuE41j/NMznhPlQZXMoSaR6rSTqFOWBYaGbdiAL5RbneT5ifQS5DH3AAFu97
CFmc2y7CqLrfvIt3nALxGm1fcGd2q7w2JbYRKmscfn6PUmL7zOrlY0lpTuTqV3fsLmpUn7AFlrVZ
+DEjdV8Cutb7WgUGLFx6pl4VqD0qPJDZ3WZ/t29eJDTvzD98Zj2MsPXYUvLnEA4qbCTKmBAabnVe
8pWuSr1VtzTkr6qhMBkrdjQJmT02iyWszQrMqb+iN7G7qkLID2OSMy3A0Xe6jlNsyIuNYcEkvOBR
a/E401MXqVen1ZluvB/Y8Z6pMzcFmtZHUmYa/pK8yq5/3eMPFLUmiGqIZEqpR9JVP4OWnJs1Wvm+
FEGXxWejnN7uoBn6Vj3oMk+nRFxolmyMeDnXCw75ObKsJXgRr/ClmsB0+hp5Bvv1Hz4TU/POePRt
IJxZP7q07A8pp0oGuULyBvnT+F+3HXrKXjekBlGgO408QTPa/F5TWB+EJX00BGAgR2yuHPUanGbu
svH6ZLfb2mQ2kpo4PI9Uy+JB6jtdlQJvv5ojxqfqPedIdIoG/jVmbHQu6cgIem0PS68DSDMkNDPv
p/sXu5VG+bBRvw0oH9lnuXSOg63WPdtnx2FVSrmXsEc2llTHWPn85WNMM/5TLyKuY0WKmu32Z5WO
uQ1KtOvKHOERXAlw3Po9sWD608UXggxIssotleAg6AC8nzLVco+tUy9PFdyVymiiIBYT0LjE7b10
BJRqtYdm8djlJOutFmesF1Ntrc8o5/AuM6o7yHyTEVtIRU537N+c1He4gBYkf1zXodiaq4hRpG/q
PKEsV1C+/Q0ymrsGtP6oIf1aH+RnOOk5ewUKIThmsNVt9/1BFerpJbAO5AaLrcn+Cp73H89Jclks
8GREJwHYqBN009jeNzCsnOnICNUna6yzVp8FVj/qFOfVIiGbN9Lcc1CnErXrdsii3snaAJYkfxYy
nn8V7UppNifgIjBFdNew11lW/vVHGXrvlZxCE2xirYDbfjU0Rk31XCbikpbnXbhatnEiydK3TiNk
pWKFJIL7SwfzesIeehxGFgQGifncjZ3venDMtfd7As0mBnhFfcFSkCrZ+2gfM3EreFL5hj2h/hb2
yslBUeWyG6PBkHwP7OGeh06LWl4PgxW2K2kYGIaIhgkrQyp9XkEMiRBNrzM9f0s5KHTA9g8pvgHj
ccDA69TN3OFbQi58qNTzYgCfE6W6o8aggSZi5MnmkZI/hBW19DTmm6z4SBS5ODqqhfmRh1f4H+bp
KHvl8ybil/ciPl4b0yfU7tsPTNEzG0TKEOA3ARvgfiOwqOWEesaoDpQi5vKikh0yPDW+b3ZFBLWD
4Aoit2xHI3/KP2lkK29TYFKH3mEXz3JJJMVDWLcf9BFSa3d0IfU0gD5rMM8bMJcnX8KwHGElXZ8b
vBQ1Ztont6VHwPZ6CXTWxHznDDX6v9IpEqyn0r89vDqe7k23myNFKlT38rOhdjDkLzQ+1fltKzeE
cBdpbtFqulsbWWoDzZG1qT7JeKGuf42GKzsg9THE81+CJ1RYlgyfLJvJB/Ox8lAFsfpm7HLciFpf
iw+UqBOKX6D8GOYjq4h6o00RlklZjDaogkYQK2j2Gr9mmakZMIJQDIGooAHemHw8SUeLnmE5s+Vu
e1k6LGBJJU8jQnWdTeeZbURkUlVNMQVW7lw1AQLi0VA9+juQjyC94eR7UlU3Ou8a574lsI33LgGl
kjUfki469ExRSZ4TygVYXQ6LMYMu4mvacKHbRny/weVnQF+G2I3Mh+2ZUiFQ+I+Xa39ftDyMfyEH
SA1FA2ok4zfsG1ue7HPAyDKgkOdr4HPS50k7PzSLpZ4MhdWkscQNK3Y42wbCqzUpOwKO1oB6/QUp
Sc/hXnfsmnbsyXwlgm9SMQ9Vmqiy6Z9kQ//6FaSAt5Tfyi6nAkTJ2WqkE1L6kVLrYnZcV8+TN4VI
UwfwCZf+1EO7Yf7aH6aeW/Bzn9TDOc2VKynINr2KY9EyzPwx0oknEVWO5IJv+3Pt3bBOc8wYIbVf
g0joo+Ip9gyGwyI6V9zY6uIn92lE04BAVSKTjUBpQZnkrl3GGiutKauMOra/xc+Iej4Z/WT2Qgg3
9tzvqZrCHS29YnXeyBUUeD1cLu84BiLmPyECb6L9daEYViKiBcr9ubdteqdsixTsKPZwuHr9I/CB
bppzntn4lN/qyWgNTqS9jR911hNjup6gHwnzst36LVfYA/3OT9QKxLRlvhmroa11LO9gOyr85OAb
H74x8hZhUc33fIEGm1ZN9XSfhS6Tsa0sDR3g5cZ57/o0IoowEaTAV4LYXUyVeEFohHtOAB6FVhsX
cWp8LVsJDS3B5OmmFQX54M2Z+f82h4yrkVgGWdbj3d3iASentSR35gpYXsENpqQM7I8jrSQ02CVn
r+z/Gno3+Y9mapB1Aw9APX5T3KK1qWEZaN5aueVmfqVj6ZZr9drh1yHqbV1sCmaUj2AfU9n8t+RJ
cwFa0+7zxpxw249/pE/oXaNb9Tisbal4ThhiPVvFh3K9vp7RaWPYXN9IbLGfcQwynxKZsJ61X6HI
MvlocK0a04RbcjXo2mx3uzjZzSefzEZyUJhJTPrW1tuGbPcZqKDrL0pYVjN2u2BkMeqBl0QxLQUG
h9GZBVVcADh6WXLgsGk4DU4szUmUOK+7hKWp6r0FV/Qe2F1zC2/xUNXeQbratVL3K1hmNtvOg+sb
XU5rwFsaBU/zpM6EHSbSvYsk/uJQy2hnfc30skSAqDbi1H/Jk372z/nAPiHb20VbDn0HCfzsZpx7
/xp00Ru3UIkBPGqtELIX1hgWyThAaHZxScMSAHPAuCdmJpN1UVfLo53wcrx+vdSZlSqLTFAkhxuB
zE1Rax2oC09fdvrSnasGsy5bLrEYBD+JMF4m4FBe1+Zf+YrXc6gOr0mQ8AoQDlmS8UjoGchp60GN
OeNJLYyUWFBmGBojNeKcQ6RXMgMzdwfZfnhIjpSRNPhkQZ6Uznq8EMa+5s34InIsCAOeadMD1J03
zTKHensmt8oMdGSHSGFrw+dCfb0u1qI+bZHlrib52Sjp8y7EFJ6I62DYU3nXNz/HYEQv72sjgJpi
dqQBnV4RTbpZxcEerjHplor6R0Z7g6Nmi0+MdFRJA/j/yjSrOEmEqtePGqi8Qef/dPU0A8ZxbiOZ
VJ3dV98A8a0ONaJTDK52m8TzfRgCHGKFmbZeP/O5WcyUZN57xRq0klWcpQ+k9GFaL/3iuCRNf7LI
WF+/9RNM0UNvQ4mXBty+6WCQFggkoERn0IY76h72LE78w3PvHjyEJLkZXCLyek+M3tHxdeTTbo0r
KNoi4vzmYZlvLIHtVZR/oRR2et+6B0AnpwLJct3xNcMGf08q6gZWXXqgGHvM0qcy4F77aKcAvKmn
fLZJKu6asrPG2+ppVzm6VxbJaT+3IGojL6iISr43336T/vGbnDwlnuMAx3DHysrBtAPgx6igVYK7
jikcOBRHmeoGk25wqYO3a/0xxSJfnz01xJTKm5aZnezgBHFh4tmc/QbYXKc3PB18AXMFujGejjxP
MWOFvdj8l4zz0hPnn4PAd+s2ixDmo2hYyAjhYpuITS4bA1syX7wmRDaWSMXnMK23HW764D3fhUTe
HqeNiOkLHK7/+c8zJG2+dsfjdJ6aI6LcOphQVf1cMNGjoHjgWjwqw7mP8pDa9L3AxrpdGWtt7Kcd
o1CRAWOcQ9Jfzt/IyF65c+ZSmi92zj8G6y9Yt/zsiX/B5gwvg9k0rYyEbYuL/vix4GWPkWM5I7KT
LO5TRUJCB/Qm2T6y6yh8ngbDoPj4jjiBWJ8YiZwHoi0+EXUT5WKRGCD6kag2O/uZFtQh0GBPzooe
x0BuCzlp0SitClHQKO6L4jskCMM0zsRJkyd6qLgSo5rbIT07BEXqTtCwJuGxdgHu+R2KQcOLRzhs
bBgumkK/Wb9K/MdqHNSmTe27aEpeojfg7Ef6x6h/cwoOv21I3Rn/D0R6+NY1EBp2XkpWhTAdLuJu
smbDUdpFDhnC8kDNaFt/n76FdFZcn4Fu7dD2WMTUyfa5GEQ22xaquYtu4kWqUZq8hyLj7HSNROIQ
j5JHSgmhyCZ5cJ5aMqD2WrexhKCpbSpib82JquJgkDXbgE9oHk0ccomnVbTIoJgCh03pt6GlBxnq
2WB1eEjDzuDUx7qhQWKEyJRXHXozUXgDCxRN/gjEL3gzGM4HHJqgj8Lh5TsuetRE8Leae8+L3c33
tFbCj/7s0l1vuxtXYV9LlzY0AXUdvzxcuUxdh1cVTyu9DFJk1mTfZOCoPZaZ20bLRVT/oVqFAe/8
XXjn0pnQ7WQK37aswL4xJ4v+UA6e0EuwJCwhTH3xMRfLr26qaVIlxmrNwMY/lxyN6eNOkU4HcA7+
KlNuikBwVK7HHLiP3Zf2m8UEU5+VwswIGQAuQ9Q5vQTNBA0V4kSVtfJPJFTIELQLuKcPx7jdWkZ3
JOnf05+QqVjDq/C7PfnCz5drSTA0MlmkoKzGDEkg070j7GQ+xgHER6dszN85kC6kmWTCpBBZND8f
o81NbbbYs97n+wo4suigQdp/ArUc0iu3WuMAtOpWNaAJs6yvUySIgrayv8hs/Yn86P5jm/VIdHVM
RprMd9XKM7jcbXb5CcH/EJR94lIAH8ktIGD+HWr1x28UcsHGfvvn9XThwyAs8YsAH3uQOVSXLtyo
GZI4vXMJkTajYMAL6k2tEaV7rgDWD0A7lYlA5A0Fc/kmvtXGACqdcxPQeR5qqOf7jTvNB6/2lkSC
CTdgeJk/WegGjM0Lt731o1G5rzFV01LWRljRetvN51XZI9ivJMq4HCiIpopMWdckh5JeZBws11+n
JVVdIljuPTC2Ju3iKkc8W1jddanOT1x4MbZ1QCzEwS3OG/JMBG9wMpwD+n1NSv3jUH/fhDlWCv+K
TW7iYf34ZX7J4rpYn+6Raq1oquLnHMyrk8BfFnerr7tHLvQvbNsQ3k2K64SA0BBo4mML/ioU2/Fn
03cB00OBb7lE76DEDBp8/nF5PYOXyuQ1tO7EtYWUlRE00kMIRBxG9fjsi4jL4Z+hbCoGOVADL6gr
1dKIjPsKAHlgocZAmaeKlh7wsdnCv1OUJObRrdJnPTTyn40CeL97Srp+b2dqDGpqT5qgxaANOtUW
2qiRwMhH4Zey8oaCs9mNOTtTOOuiAPjgiajNfgoVu12JFqef+ovkmRAXlPlYJG+lHGMzQjgVZ86G
jUsyB/mrtxklL1/7KbgfUOwYdE2ZwDrOpMluOR/Bl9qzrABr8PF2pedNZb6ctXvzuMx+da7mEYP0
AInmYS9DsiXiljUh7TSlfA8dRqFonamS+IM0WzJcgJvMMDHCVD/F0j+lfVmqxMtGuW5vaPxGaRVo
MFwqgnYKIP7PhXv5ccgRNY9xc6TaUiwG4oq7NFP9pdDVUqKjVDU186BblubpV9GaQl6WHa0YEOpb
QPmkicPb4fGgyBoESbyR8WetaqD9zrUpIGGhlvYYQ8fDHT9F0NRjEyRgI/Mm8ayKSSReMZJoCqVr
c0HQ+lZ23JP7ewWkVAm+/miib9X5XlqOm6TWoZpvNYsLn12DXGnkFcD2Kw7L6xA3vUEGjPkZvmfP
5x9W8qhoNmHpXuQMSGvds1MJdq3xbJW8+W0rYTMw4STfbR1g7uceV0sbZCFNPdna5gzg8I+njUzF
/NpJq/ckNG2Iz/zKjQInWvsoC9hqoccKHInioWF/urb49+s7h3CQSQBthyfS1hr8aOs7dvA/bMdh
gaG2yPwIme3TfysTtVOyQwGG1NbPiCRxLRuU25iS4jxjCdDgTJRhZ6YeutlKjjz0/4oB9DEikhaM
HqGCM+2katXiiMUwMG1QSoHZmXRSAlvvu9UzuPiaJPSLOHBa81o8ZKm1UGVgfjMorbPJ2f/gIJUO
4gZKoGqJYFLwYRMcEDVl8gf0MMogx+ghmljR2t88G5osA23sQFevXLsoNWSrFSBIGUEinko061kc
z3pP0GbXh0iCW1WTLoRepBnFMR/6pWmw8bh52/rbF59pGD6qTzIA5fwmmVfls+efbHitP7M/6lIb
A4e2AKkeLuuYWvr/zMqTg5lSTU/t5CHtHLaESjsCNE8pB42AdkrxH8z2FglCU74jexVzrKOCS4tt
uRI0ICzkBEwKCQzso2lIG2UuAVSHAiANojYKf9iMkYIneW9+0jpHCh+DpdvVm2thfUwnWZjpmtqy
+NePNrForLJYJGfKBfkNyF5ctOHZhLkjqVGc3/HWdufq0PTaEIX5xfRMsczVyzXLY9s2rGd77zMU
nBNdPaC7aOEtsuEfKPDwlhhRtarGo9F7Yw557vq3irJqptUfU/ZVlxik88bXXhIL16+o+bCc9boA
JD+eA6lT/SDZUsN0NjHEG00Tr/suQYTJe70Ztaofo100pKt6XjRRQIhHXB2MmLfo3eR6igjdHC+f
hoYmVR9MXTUN0RjUsaLdAnv+pGTtXTWHdAX6TNujlVovzsRD3qjI3/tpW5Y49XYALAx60Qlvnjz7
zmE6xkSnZt6oh4NF4Zs2dfyIwfPZ8V3dnqLFdIJjgg9Hd3Tl4VI3b0qTP0eQ4rPI+JDKONqcHfiP
8Oq9DLYENWCGTE1a7vU99TqQI1v7PPWgQMB8Nbl6cj2KaI4/fBCGkVEDycO/+iOLT6sNFNEcLtBO
dIBA8N6QSY9ObanySgJ0ITxeCkNsOZXCGXeGRUoa3YJYuuwK1JQzbDi+J9g9NAGNf42u6DAriOsO
dx6sr71E7MxQDdZh95TUFEfvQnReRptEAwQOGgsvmhjh5SwxjGOsy4kYofHwRnfE+OCvYYiuJazu
6INKW5IyTpzhoApxgyRDtKud2R8RU5ZWyKlT92Kdw9BYY3TRP3dlTlJFUxRdf/by9RgWDQi/uGJ4
Cf+i42K8wIPPHxm6ZFjaaTwOh9p04B2QTeswLiWmXUFoKo0EC3USHPJVnzlYeRHxpNhmur7rJwET
Bh5hh7VCurYRe+FMJtr1zvINIzMSpBt/Ynn87ehsrL0oKODwySTZ1NiLnBE85SbPjuNa82xEh7pj
Dsw1sHwxF6M6Xbwn9NnlveazLfmKTjovJFRuI5uSx654bEB4wf25JnqN8DjbBzbWpGNW2oPjNKc0
DE0ibF2lycXGoB3FyDmzgq0G/oz4x910qnef6XnCPixk8Hw7tMcFTvhKrfUBhvggA01opmPujSzd
s9ykHAG1r9kvggUiQexTYXxjJFG4oGP/njjjoKmkSAIqJEOBvh21X00L4YEEhwpFEqgVft0zXlLY
mvKcdxwp1nVG9VQotKRR4ylKQemZP8HT2vUnXwGWS2H8CCAdNIsBkZbCmV9adixK/7xJX7FKy+7v
Zjxm7q2O8ZNVlrCaY0fq/QRULSLpeHzHUokNoZ1nRNwJ+azHTupgiHz71H+q4kFOiifmGr5zBroD
NmD9TEYxDeyESuKK8rdZZRZ77etQuZ+gILTJ9vukAMO3QS73EOFDW3OMPSQNvK98XEqoav/IHvpe
/xIaZVfVxkoVgKvd0rPk/OROdOTltFq1msyLAGgBFvaC+HLAJSOn3zTUa/4oc2C3jcINjqAVFOV5
8mBPSVfsbUHRF8/Ygl8lcZtKWI2RazahsBq2TcvsZRLMlzYbsX6xtikNgL6PFHQwn8OYcG5NzLtc
/hbaIVX1poXwen+py8POSBQO/J6gvI0LC5CRnQfScIsb5MSnXSa8gtBvRzcqwYhsqdyz8zCs8aWb
QK+ss9EFrcaCAiVL5BLUJRbeQnjFAoJ/uweYtDpor9iHhekrDw1YmDYVNcK/CRaC+B0H7kObxodf
0AuvRRDBO2wvjhnV6otu+sCLezqOjnOMpZahr+MAYm7DZu+GkxRMJhIqdqPOry+TulMw0uSRnoLc
oepdB9AGUeTF7M8+rE9BPb2dXFXEk7AyNLkYdhIezhOLMS/I+ItLRN0OJHePc8AglRBG1xO7tR79
ki9B1eBWi3f7B80KodizbKfdRcPsvJ7+SFsEK7NoAEtqq5Q/C3u+SlERf7GfvTCqIW9BmZcb4MDV
oAAEnWWJYA1mMio4iOS+yGShPV94R3J4TLrbNEy14bZmFIPEoO8s+8YwZDz3rXCLDNJqOOMtKF3p
qE1YX/3mm/ggtcq/i5yXfeTDjLfoPXsMp+y5hXuvmhkAH+L2onQy+tdQKhNTT3enMnDRl96IHYZK
k8Jfh6C0gi/bfIMoGKllEDTM+ymd4hHWRPhk/EP/WfPwesMY9hq0Wxrgpd3qew3dv9yarRT/sdCO
fBtN0MleiCFFbED//+thZSNrj0BJdsevWtXh+5iP4S+URjjgVHxNTTj3Ue7JEMPTTcsNJk0Qk0uY
ZSn3UTYrQPwvLJEQeFWABdKUOtFgo+iaSJVD/DalAfHsfshMP0pCG/Hk509+AVc0nWOksMB6vUtP
qF3pMwq7AM4XD2zbZJeowzh/fZAMbrtetHD3apbQ/kSrXqWHPUGKmKMd2ahuboyZrf0zVOHwD3z/
NLIZ0KDbWdfNikixeM0elst0067uWZzv5XxKZDUmlhZC+mKmXGunDSVffvpU7Qy6YHM+H4Nx9eEr
v0136HANWSRHdKJoANh3OjnBYrtKlHf+RvFqCw3BHpChdtZ8lgp411oXX3bEcIptJkMKmJsHwslV
PJIaa6zVWlFmQTRb2oQYFaZMgpayaVYQXUV/BKOqD1v+3DYs2GSVUaHHS/23eYA0RyTZB8l8v9jq
wBkiTE9dpkv4d8R9+k6be6qUFahG1Z0zYfbuucUiORAtSRUf8YadjVub/Tk0jmy2bpUF4i9Pivfr
YE9YQqQzbclAW4huuW+kqICBiABeFuDHFFMTmwvvwp3J9mT8MOcI62L9LiPUHfKPEz0zALX6A7aG
Mth78XSMbPh7SX5UD8NOS4L4/lISmym7klmAkp2W3Gfg5H08Rbt4X+ReiHcqNVpZLZOEDNj/r19W
6I8TjiffmoAvC8OtnBcNdAHuR+griormRU4uEovBhehWiN8p7NX+NeKOYuf3YapjdW4s6qMH3njy
BmU4CzEs5hupzjMzuTw3rJ6WtIaFd9Gzg8/mFBuh9TFnYaySF6KlCXZ4644i1WAdwFfJe5h+tQhS
6lRsetqBJ3yrQxXxkPcbs6OdpoKKK/DfASoDYePKszZDSo8Yhl4o48iiv0aqDAs8tBavGQGFl9pK
ixSn/NxztFXHZm1gXKJl4S3hN5s8P+fTBNJ0bC/DR+RATZBGg19Qj4VX+KH9YbfPPmeKuFTAkzMO
M//Yna/IhuIaIhn32JiMOlm38yP25SInbHcJZLd2FJU3K1qws4CZPZkpGmD/Rrku8gu3oLPt5i6T
5qi/bvHaHiyz42xZN7rCQPCW2dcf4ju/Ih6Ragbq4SpTYUJbiwFeEu0kjP6+ugkk0+XA5JeRIP15
JsPIi5mTnDjldu3UKvkAiLnLSt+FTcRaW3ErC2KbLC8VjTKEqX3OB76fqIivbIIL421My2FPNCbM
RzqUFytISxq34GsUbRDJ54YISfcmNbUPS5U9SuygEu7Bg9kR7WBXOxYcfj+qOtktpYggxHxnykFC
CjA92vauAmHgZwGAq90fYININZ3F87WMUBEjceBZHzV6Iz2LXjztcu2XP6iQ5j3d9c1QoXiAKr+r
aaf6qAJM3DYqLgLtRE6yGMFuSXsGwwVVCNh2gW7eZE2ytPQNfJf7+FsBZUQci/q+GzfBxLwTfbOA
Hl0H1NqtZLkIXppVrgW+1xOXTk5LkC1L7jJEQfKPpHNMiEBgS6WhfiD35nSVuV73VATBpnxZ4mH8
ze+Lbsptbii6hIO02IdpajnmPK5XlmlzCiR/dBFYFbS3eq6lK27mGRVSsE7I/yrvrR8trRrpy3+V
yn9QwDlqgKU9lcLlI97pkasS7rosdAcGfyUIjFejN4/8p6wR6fXxQDi3r7NBVSf+Ch2VedyYQawd
hiZVnZHRI+Fa2NJuqeAuY8uoisFveejxgUYXKgW6tta1Z4HPFGVix6WhKnHdLhSQnC1zbhRHF3Pr
BQbSxdCYdemRz3zXDHD6zVCw/mtquRNLClGKnt91ibjScgh/myvOxXZjsPIIb9sCet/6JMfc82Lz
mXaE9rX9ZANRSRRqMi/fwmsirPt2ktGX1KMs/YBQYbIsdXXFZrAfcartGIqTQQJ4d3J8WhWrJQZE
JYIuollBo//c3b3okWCocfl1+kEmjwt3s3Qhc25XdaUncTHe9SQ4HXfd0+66aKZo6hJaKibRq1e0
uvtlLoDPeF3a+IYZKbSHePeu6WaUUWIZ1eWDjeE7kpQ+rIwaGxDH0StGCA6XcnqNR+xpeydr2h6p
gKfhM/Fyy+kZo0HyWmaOj7A15k6IPDvF2BQ/U4IXJVXdeo5OLym07OX8HrNAJErA8TAxrpbSyTWW
tjfZyRN+TdrWpCf4Qih5rNWYtrGRS1Drfc+ihxkLd2gtUuuEbx0M5jzCJQpEH28mbHXG75EtCtQf
S/I1IHOVgsp72SFtq6NteDpoVEOJ7lucW3haU87G9KaFvecJwVsrkxLjyAtsDqC7km7JogcVUz7v
mcwuoF2/lKyo+6AdotYSjTlxqM7i7izRwO0OBuMQjk59FXsqNrLJ7qgzQIX4HFwBYiwVG+dGnS+3
NPczUR5FvToh5EbwlmsCM1lmKJZXoi2EZJrGlu4Ja2ByCSaxOuAmhnTaINCh5H4OuG12i9QbLmJ4
ataz5XxmGD/jpCB4v29E2XsLFEQWPoRztPr20Mt4c1PuiQ8SFcM80UzdwZA2uZ/xq2rX09OX/kkp
1NgbYo2FlRfJj6UKDxG9VlIkpPEX60Jxz5jEIc9xl3yGX0mFe+sN/RUyNNqT8DAx8Yf034uPyBw8
YQtPKOfUsBheHHKiAnQLZ7eDy4JoH/4X3oBJ2FhD483mknreWg1fVXWx3lthabD3+q92Zko8fJpS
/csXz9mB0O77jRlTwW+CIMd7Io01b6dQz/0qx0oKG/WS+m4K4TyWKf84K/5pmwutETEiMFCz/vqC
qheOiq6AxybMfXh/ZDpYrer/7+NX/gXodqDZpk+4hOrlQKrMM6NB8aDxKjeWucS/n2VWBXEaogu/
DP+xj8fVk/xkLGbsUQmeDxMgOVJlx8hMXsjQ65a/l91jMYNlNKjMYFvJTu70q2vGOrLx1xDHnDsd
foMIQOU2cBqQQhDS8WReiGo3a+ctWIhxxWtFK/+VWIyX4phXO47GHr4cOEDjgo3u/wI7YAPar2nq
Pvk/LNt2nDydA0peF50b36Nx02lB4g/Xx6liVAYPullRlnlHq9etuUS2OMRfBWZsjhR+n/W0nXEI
uGUeNSmAQ8LVtEIMhEvlBnwFTt6zljF3hUXmoq59kkY1S5bVf6gcJBs7PFRiwjYc9JW/IOlhvjR4
42FyNaGBL3MVYP5+Q5Od8tqcXgBU2hjab7MWfcNOoRM4yH0gdUIkTSX560kCZYHKqrV9B5/n6gAU
IzOiCVfRq0hjiaPVSDJbv1Akxu3cZgUI8LlVWjUJoPfO9l6mqFrw5HDATXW/NT3PZ+mbne/y/30/
VihWbzhTORUnzYK3l4/Dqj+QlBv9OEoveAgH+WD+hlWca1GoNPTPykiK/Kmus2iVr4FmYPQ5NfEO
BQYLRgQHnpN7CPDkIuk2G18d//sfZJ5Pa3O00RC3TUAQdynIKTpwF3bz5LDNokwu8izOTFmFGxFA
uOx3BLKKHPkzHUXAHxLhEbvCb4C6n2AWwkoI3HWTbm0GasO8dQ8Y7wzz37n7QUH1Dv6HA1UwBgw/
rZst/hK3CCmA1zjVSut4eXlMbzp7gGOAK7sloLmGozwUyTnpWAEmrPxmK/OwHmX9QgUTsB17frJw
BihNu1Sgyx+rWQHZ57GNRBeqJ2nZSabuyHlXgq32dERRWv7QwtYB7mTZMb/cqh3Pbw8ewxdQqARO
iq5RxGH0A0rhrUnJ4vwVfxyo1yrczJ9bL0kyaoKECKe9q+zf9rhRMWbWwQKi1Ds88b/oBJsBYj9j
/V9gMOUK6uDc3+AtpFhAjogERpMxa2dTIAIGwiMHN5XflZilt0cX16o8WT2rxPa+WGxURwWogGBr
46wEuM5iDx5+f+pWJAFEYLd/faYnkV/4DXXatOyiPkeOFoVDT9sj2fVNxermibDP6jGGWqPWMjyZ
qeqAMk2UCd0w/FkkkJDzFXAPDwACWWqtn2TS9QJjwt8m8qJwG204ukqy+3WgZz9h3jtCS1OjtyOG
j8jO/iJh0I39LG8OTlTzL79/FqasArxQZjRLLikCEMrw1y18ABC/8jpCmz+nHFxkkRh/PQJXa+dW
QkvqPXW2KONv+J4Uh1aDgGyOoY88AW/jXcvYJOTA/VVMgEpZgpvnqUzHLlCI6kKyI1Pb9klaEUcV
It4zcr2DOXIRCO5GpA0pr5enh4ax56I8xEfVpw8mhNBhL+yhv8iNNGormEMlWh7aySm0zWLwV7Y/
qKM6Vf8NyyFeRpcs0FJHeynHWZod7Xql8P/uKqXw1/TPY7g90k0TjOjxeddDC311O2sUA+YVCswD
0Z8QWxAHae2Iv8CNnFVikxd2GIVEPybJNEB8LSm2jeGl6hdJ2Bh6oGg+XuYv7J+NTegHtt4RA+1g
hjvm6RiTOWA/+qh6zRdFd1/LGFXF4r1vfu845jc7OvmXu28hnCO5PwK8gTVonzOOWkwwwg7zb4S8
tQHEcFGnRrZg9LgVT1RImLJJmNNZI/6bpsWz5BysYg32ZEZgBhX+eThLFFE1uFz3CaEkVCrqHZcu
Bfv2Y5Dki/KJeuMrFDgCneA92k72DF80FtPAnlKDQfB6gc5ub+hMUzUkokW47rjnSckSJjinvtjw
4/qBnm/42f0+BidJ8PVlKHnoHWWg2CMeWyTIzfK9aQFaRy6DPmSSVH8Tt5V/FODOue7hdtWdvqzY
YsP4skPJpiZ/B1gVKS0yDCxg+iW6Ws/pKDs8UFmN9S3d6PavmmrLY+N7ENMaexo1YsHf+KzLVOIy
YjsCpFZ+FdHcLhLbJlfzyGje37+wV28ihDH/vw+nGXdowss5YHbaThQvPBESScp0huz3D6SsUDb4
NcNpX46PKMffpUevPgDhJjgKaOSdh34E4ou9HpJOgHUZhktw6LKOVt0/L+nIZXQNIKnEwomxPsYt
ZApko3is2yAL+XJ4ZITcXVv5BYjk0LrdEVHH4kiGVE+iL3UdTEnoQO8M6hgckR4j/5pJqby/ZRQt
dNRsRxlDAza0QJJ06bRDZgK8dI+gisZIVTnRVoblW8h11Kkd69wb2Dpf88AnEFUrjJ3PLaMYWbG1
H8P1NArhPlDlt6qzte1KAr4lArMJbupyBOgxXnWjVqjH2WfzqnrrsR+LC5MydcmFASibZlufs/K7
75eI7ASrt+30GxRN7u/n7a4z1yFNmzzw0OfuhbCkxhEBi7o0XHVVacgOLzGyRm61SBgg2ulC49U9
1D/FLOgBwHdRQfaiu/HdZKPSTIZXo9KJ8VcRm5NRwF72YCH18UgZRK2vJnpvaEToyppZdT4sZFXo
pEdk0hxIv8psmUZ+h0VNmXL+juCpjSzD9ttUtO3GTRms+KJITA8DsFM/OFddt/UF+An+BJWJ0bqp
LzxWjZ4tsWwppua6IK4zHxK3pKFo5oIME270KAj2jYdFUZ9BOtl5CSSz2V/pG9uYS8Y15cU1tqaa
TNbJ8OHHUNPao82jeGS/gDKHY/mJa8vm0UgZcPWnBQr9lj+2uFPFMcqT1w7QznZUTs8UH+z8Qnay
PSa8ydFRaKSlT1RdZC1xjzfhf8V6zpTjXfYHCH7nLtMTVLYtHsTw4Rgr6uPbQSUYzpcBlQC6mvne
7oohUyE1IXX38K08tNaFbkmvt+k6CwjCmmkyjKbDR9JT+BstRSFDlIAOM2EmcRp8P2IrQNEd1xgS
StBiX9HxbDXBbYS4pdHmpXUEUN3ET7PlngNKRy3qQkm+IZPRbo6LyPXKAg/RAKRueqchox88cE9e
lt6dgNbDX2BXFd49mIZOXFEdx7EbA5xOd8QQVHzjwqoWHmasWvt4U59SbpLUWcP1sjUFI65gxLY6
R4qn7UQLVuNDinH6lKDNTliSkgeUUGM1OuC0qraZuWd+zlWbLfNqpq9tZRLr745weeZ81oF8iREp
gfanfxMC2cqRE++ysjo99SpUWzlgQC5kZyRzliEAyjtlAolXYl0vqeuFbI2hTPtHpWu9zSFbOXyA
raI7Ig9p13+yX7sEN0+QADLsH+VAuUEzdSMDvjgZSUeQFoNuRxYTJojtJpVDwNTLdiQBlE04RhLh
Wm/qCBvjj9ZgIiankwq/y3dSYOEQbt1r+7pxySj3cLgXgdAI6iLnosNcM9JRUta1b1KwSvwpsTzG
8Xh7jNY5NYHo3b9/jfVETRL3+iUlhlWFhj9gg1l6Wia5AI7N1i+Cu2aOjt2DP3pzTuLG5ktiJ9ZS
ySkjtNRps+JYujjm1hU5KmSa85bNqRrmO7Q/ZPH7vl/QGtdzY3mjQ5+wYJMrJpI6FWrb59yquSUo
WkJiDCk9DzZIVvS7dhGM87e3qCsZ6YpyPQqko6DPFDKGEr/zQPikp1Hm5WxLtOWPcRSQjB9QlT87
7Jn832V7NyRGA4x8kV4FAM+znXneshD2LS1Tcv7L0XgoRiSljxtqT6RrMmtN5wrrZBEghY1vj8lp
zX5lieNE31Bi5+NF6cpr1/V3spw9BUWU89ufAYJ8F/ghBZ9s1EckiT3pugaROjEgH90UsU09+n/J
LdtIbcbG+y1SXVD6G9m18G1AU/W9V2aZUKk3JnnGQVsYT6j83WXpMxYHjeckOMutrYWooUzKJT4J
12F/4YpdnhGctDf3ZK1cXsjqOCtN0eL189Uk4PzR5JwS7DLK4iMtx9kIoqZcOsx1Pi3elCc0z4sZ
c7bJLuFsPiXW66duDYVKddNV91+q3pG6shUD4F+lq7HNYdb/61TS8S9MwGYc6gyM2bH0Q/1vuSFz
5gv1wOmDgJFXBL9GH64C1MCbFZtR8EGI6knEXrMNqIvJFRxKWpUXC8fAMUjKz025Fcir0IzkzYsD
CJcHr1Plh26iLyHUeof+TwdInbi1FWPR4cs7t0CVH/8vKtN4w+PuGHh6UTKQ8PN8Hb5WkPR+p7aE
5JoOt/eQEHJX4H1RctetM8dtvXfbN+noBy48gJqzkkty9VhlUaTrC6c4SYbas1qBjOiBow6GmY7e
0XBNF3FqtklvY652cvcJfQstlJdFbLExUsJ+klCquDdueCtEQprAFq8Jqo56LFwSC1Y+fIqR1wxE
990klIEOWeluTgQIQ4Q75zQMZ2GWaNkR1cG5AhMQ7EQLdqjNUS1eWFRINKeq6yktc3OZ/65nSVay
M7w0m8khcABXuihWYlTx71j6bKUh5LO0lum75oiSwscAITg0jYah4eb8pAm9YmdLydv7td5PI//B
419FWjnhEk5VXR7NEYFmbp0pLHurXaHsL67MSrJBXr4YCRq4zQxxRnha8MB273eZpjBs07z6E1vB
txlCf2KmLNd6sA/ERAa7mLO2zs0g8Y39azvmOVpUtjVWtWsXTcmiNtFFgCVbll1/4Q/fbA99iitB
CVbXo2jPKFUB70kPsdFpMIiFmOlo25BAYq0x6fXxMUwZw7ywy19cvkKXMS9vERlJMt4b2gigJU8H
XUVqLAE4vYfQKR9I02gt/vSukfZNZ9z+YF6Gqk8rhBrgVJWN8kV5U/ASWnpiyLvlv2nJpzior73D
6QXrwAGCFwbR7PiO6SRHFHOlV7ElkS+0f8Qelic/ou31aUC1b445EGXm+l5Yl7QLoISvHXPAjfx9
22Bv6sLZBpcYxot93LZotb+Bc665awZuZ3ZE1E5AyDL1xdgoZyS6azeU9Ua9WJxGflXVE5zg3ANr
Gc5r7vUbA3vWIvPntTKSLkgSuQGLiKFDpNpD1sksjniUA020nM8qBVOTupbwpklxfAqAA24ZmNSK
OvAbl2cpiPwbXGl0u1qMj4aKgggv2LGGvaT/b9p6qdEC4eVqE+UK1cxCXVEIWpjqYK00Bh5sJXwU
noQ9A1UkW31wrkHQEMKBRf9D9Hoxzvmx06538dzuqMkf3vegvwlJyQe+FfXNdRHJzBJ6f7YTvySw
QqSw6VVO4bJUy7c594kEjfaJOaTqqcwyUqGgPVRBXqiUNJ+YuTkrmYIAbvGkU0npGSWpyrqIbB0N
/cCfUWkkm7yDREIgq5NHkocyBduZ1gIa6luXJTJ27Bhqx+6wLz6Ko7Smyevdo7GEsRPWk1XupZNO
1Jt2dbq3RhN8IFqW0WSoF/ra2YdmLcbgQmaDjBIFajYUCyWj4lfL4drkYZvgCbn8zhSJWLbpExuI
due2GFcBSOB9LFm7NdQ8Lr/iwYNd6dvhFMhxpqTBpb3n+Je+t3UWrxCDskWLOX2T6y7c0SJzg6We
CWtnvoTMo0uZ7+JDplilxYh468fNiCQz3RZwaDJJ63itcS8AC1XNacOvu4x61rSsdF/bFf8+k48D
R7TCVImZCLS4g3Iyn6YQ1nOSRv9Cv8zXL1nZ2FlYuPdoEn0RtJA69eVu+BgHaUWWJrKWO5oeM6He
0CGL4+Dj3hzxhp2fqJhG9prvDL3yZ0jdhpXiLzS9QFegIgj8h+mwZsOy1OmTnDwzIl910jIio7ID
f1Ik2xnSCZ1wONJ4/NyJ9582Dp3SCGL6vq0LCqGPhUIrb2GSYElBUgpIV1ze+7InFptoClfZTSu1
LlktLZ1NiOsu7eqUaV0cNrC+0uDvEpXRdIN3qU+KrE3nbtwCVwQfmL8BiR5QnFGr9yYyQdW6wxel
Me6zemIZVrE7jtFAml9Ckak43vl801rJ/Xkkt6BT+qs7QkhPlOJc31JLvH/Z1/ODmKLDfej/sRXA
5JcBXi1dKUg1nSWsmAWbH2/IqvvLM6bGZAC477xPKdRUclNt+55bPjnGwjFfi5IbALq5TKV0jkNf
4Td9iq9owcUev/d18tRpMh8vCGGivLRqnXdfu5kxKSUPpjUN2+Shr4I7h+yezmQa8H3h92bFarYq
FfM47VK5+ClzBPvbalTbnOPOzfr8JjaeaNgZOYkeiZTqfTBiC5HzynBvCf//bW+qsvPW80TuCoNR
53tGXEW2SDL7uO/YVjjP0Jj9HO2I6b8pseqd/p+axmPTOwqWbhcHfpWA5GNpHkiIxBhJ+RdknsAS
7ujBUfKcCItNoHNJIlV5n6Ay11/u2B1Bw/gNlXKzOUr7dQH9QHXJj9ct18Kn/p81ItuRTslahCoH
YeQxqFT9e/muy3GAag8gx1E6/p/5bXGsWqxGqiuuFfWTPiJhR0DIKu3QWDWY3111UYCj00cncwP5
hpeq8nWrWT5YC7CalnKUojYyf8mKlBLTru+KRiy0oD0lzxK3RarlaVkRXpQHVzIwr51Ob0aRU61Z
tNvEo4WZILZph85x1gI8HWyMRbCrCarzPdbYKsxi6BUjBq8gM5owA6CEm8+UOQ49iLRyTdvxNMhx
99BRpzapCQTQvujepojyU4PBkntI8WyjPAt9g5R04iz6ub3E6s+P9OJrmrCZpUIMyNsBsTaWE7Fn
KXFwJ7dFQMw0ctwe8xGbcy0Ep5XnbVrLZlktoCpiU+Jf+CNy60n/mOxOvQLox+LWRf7lGRoDMGGa
RO6T7BdllTDPnTej3tFxSjFmsQavOeoW07T/08UwxTMObeSHHFR9I+HG7bipF24ZVzXiThgnZvOx
8dJ9SdHk4WSPXswNsWSYR8iXIAuaoQjkcnlEwkA4iv5xtIjxx2pR7Bx+/8YFbtgOyKGaJrctCEbO
fiye7yiBILM6H29FFOFNyh+WYHO9y4sjsJaDZoGTANkGvdVZJwhQuXPXhrNzyibDGj1/sFbHujM0
wreY8I04BBg6QtQJxmUISXOmjYrMa0X7RbsPt7s/QAYEAfFTj6V3DN+qe99ETpjiOxyHliEfeAz5
qOJcU7UN+5QbcumqNAM/59GP3wb9vDqDUJJ5oB2kMWjQXOYLOVuszwV0KqajSR1UDgdn7intJZDk
vzL8cKKvOxAyiyrjHjUKLnWVY5rRR3N+SC8Wc8wFXAc6xUFc5sBglOwPqxh9PMQf81mJCQ0RnTeH
eKr/RHk7bpdpfkVyCSL20umqe1QaVzxg4e3RJjHytwPaoBcMUQ5jJu4f3vkvfT/FwNCCJ6xRT5Yb
3l3X/bLZE80x5bfQZDdsVEAE75v256ApLROyuuJGw65PiDN+tU5wuR7QHpgLwmPFyhzrGDgOjE2s
Ahnd1rV1Y/uLNGVK+5ZEN/jPYBIvAfIu8vsGLlg7W0AMdxCCANJ2NXmUIuP/SNSqwvMVeFf8a0YT
HjgRoKlk7xZJX8fIgCMSLaAOPOXRgK1H/fVOu32k+mGbJk1oDumkYE9VUsMUl9WodNELgJZyhOmU
4+3NLiQPY6376KKButXEkgeHPQjiAkx/A1Wx7nfXohhqnxnA3lzHB33Mw1BFTNdrhjF1uJr4lSoH
ZaMha+izxm797z2Jiw1QiidIJ9tclCvlBemR0rLzCVQaZgUaY3PVhr2Kg5RE/HHAh7AqahjBecQA
wq8akGzDp0iDlbhIYS74nf8GvMtb32p/qe6N8N/a4WbFhKhfXFv+YAqR/qzd8vlVG4JMHt7iWVAR
aMC8eZisQUlyOIG5KHppD94wt7m1pXfkYs8kUp5S6WC6ZrIY1gUI7VG0vh+qe5MvdJfvrQCvXNyI
sG/9OzVN3OF7OQr/ZTlqDIpZzYbXsPl8G1WdrlNvKKCpFSf4t6cjYf2dWUz7oWnFPdWDyj2hHZjU
F1qYmddPw+cL/aVGA1ukKp1Kfi0k8oHF7BvvTD851rM0VKJf4qte+JJS+Y0aX3EnbB6yVWskUOU3
v49tBRyQA6lCSwBY/ZedIJtttTb0FgX2DRRjZXeyEShZ8XlexzvGOsyGwW/icMeoQ1sOAxRhh1q6
2KonZKicUckDECxgKfsQ9j9/nJgL0xLx+bZusDDJYF57Nn3vET8fXnSjTrhk7CBhq8EPanMXH9Ws
jV2lKwwQ/XMkF5h64eOgofVbBITxPCtyCjqgeRPWNOWByRwgGnX04mynQOZ/r0RBabEvmo7xDsV+
FINpUlFXq6V3lhva+LZvuELfwR0V59QGl77lf3DBoqERLCf3WpaNyokVRLTSSbDD0QG3Ux+wxjMb
C1rEa//mNzt+hgFcjhRcYbfuTIyhFeU9fe2qzcVuaRML0s5bvhsvraWxH+Mn6h9k2HWqUXmeKmRz
09ORHFCPhobyQYgMqPf0MqubSHmdbk9QEuNdmdqKi0ln5DS5J3/k6QtaCi+hCV7xV/wd4aM3kyrZ
iBjb16aGwBKxYVcvhifGMRDemhEvlSj5l23R+TJ4mbTh0/SnKZOfAdtm+PskRIOEuBLqJPg+2XTf
0kvRfZghryeyMVZ9FfEwruu5AISaFLA8Qh4VT92Tip+HozgrIFMSgRsi9MuqPjHsWV8Xh3I+5APq
vX736Dkll5YyiuOd1SzyaU3+NqfTlj7vMBCRToScvQl6UVcWx+jQTAq+8Kopqux5WwTYlDDCv3Aa
74/oPn3/xHLW2Ao1uBKCm8mGAsFx8xQtwM8JXoGmXWBHztZbBujqiW5FD221mhQhAcM9DafGGzbl
CkVGUJ5GV+GjbhAEEQdWibgf6wVr1It3WTJZrmMwD0Rsex35xStZbzFqe98qPnZXz3uy6M/1sjtx
xaqyXxYgoO/edo2NYYDq5EY7CVKvcp+wMgExfPX1zYzdRzYPf0JUsyGCYJQkQKv7gRryvFKf6dxQ
Ihv75rVUdkJf6gGsBbYPEPTd0r/6lN2wze6p3GvCn3NVJtZ7X13+0PvYzpQ56NJzP0opSSg78laG
x+IQq7aeQ+2sSfXYPa+vT6wDyIaVNM66t6M/ZNI4e4VbwmhSnk+kuB5zcNP0SWyTEHz/OFb1vIGA
ocqwtEfmcF8zQim2viN61V/9b2dvZKFWfe7HBqmp+fnjJwMzq7bSQ66+n8j/Lq3Z31eeg1nRb2o3
Ur0jGnE5KPNz6HUI76Etj9v2ViXAucCLvK+MvK8a+g1nk2BORgRQ0glZR9AuAgriC0bLElgzjgz7
7kx4tuaG4c5+66NXnCyD5tKAGkvg9X7SX443gdNrUlM3EtRUe0adP3bqHx3P2HJb6CPmmOPqxf0i
EnK8NJ70c/+SjS/oPfsxUMC2TB56262pGEELL7xvd9x5L/tiMMG/W8XnnwNq5iyTncrx5HaIibik
2meA0WuHFCDpssNDho4ct6wBhYx5B/JAm9xj/bi46oV0xDpzB2AS3sDZF/cuxsDomrHZeP2qGyzO
Mhf+2gTQLNyDzCAFdMda8zffQlB0lgyqioIQoVuGXCVnTL317WQD6QF34/KTOiGMISmP8HMziNP+
i8pKfeFfXdiHqWXyvc4U9tY4Hm4U4d9qWGIRZQrCkDydl2L7ua2FvSTi3WiIqf958XxSbmLAKM51
RDHDnKWfnSR3hJps6vj7ltpYiN4sBE31n/xn+51tiJXVyYoBDUrfCSLn9tVF1EK7gDAbYPRdctaE
msnpu+V59GAWBm5uYGBiPsZ+HxxSpwFaU1hetbu/r3mceNkJszFO6OTrYvQ+76nN7F926T29nSLB
qq+gpXj97LIsrc6+BD6nHyohfSt8YeWZhkaKp3wG1zVQv4+fORKdwtFVWb0dhizmBE9u2JrFWLoo
3wX8UK+vxt56E/nnLM5VtE3IMTchMfj8Cp89bGbunAlb6shFxloVfi9gcCQW8JgsyoqDVOhRBdxK
fb5fDPyGB0LOPDGI3n/Lus16yIvRTgbaB/o6EQRaWQ4EVuvnUCSn4oPhNhPvJ6EAnAINh64HKGnL
3MQ+yuDDuGTxBUYpNTBp/L+mYAkUhW6NHfWAouINJCB++Lteyygshm8LL0PyXdZmxxlmVin+aPRS
kUZxgizVRVF2bsArHg97j42riVZvfUrMyVoATKDihDLuu4yEf2Tgz3YCCBHlM0Lw0Wh91CzC7lxR
Z6I5w/qnwqEycbDZis3etBST9RPs5wymZqDVXFApxFu6/MyW63JR7LL1sWqOIXNgH9noeqLdJ3b/
b0mXrhdBdysCgDj1bYr5GSleWao7ukZ2B98BdPLswDSlnLQyUf/Q2BzmMrLPmglRMhd5tuIyhZXZ
Tt92U+yFn6uPCbqSmdRRYY73j9AUYJpmHLnE5wqZYkabx6CDJjd2NRY3xy2bbMSEyMHi4Kk77OB+
jqegILN1dk/hbLngZU4erqaLLByqvgJa0K9oxUpJwPP9U9UjajD0/A9Nu02rPROVC9b98VI8Amvt
YSnLg48UqX1SvCgZeJe9ZLMmASUsn3Y9ZSg7Ky8vNzEOKhChEi+NprHLO+T8cQnc0n/1o0SCdIpg
3WMLntpwQ/uAXWgkm13XqIYeZ7CEC5qNXf+s2HTcrZFclws3EAdegOqe0AUbHFrjAmXuuYyIQNfX
qW/NdR2xBtNDGfkcfUjTVQKWOTFkoR2OewZkGDMuJGFt3in7KmMl/6zuCjIfGsTMZXnEpLZ618h0
2Akqann4/Ww22hAYrgN/KGA0BGWlhMXa4R/9zIwpbagFWybk8PLXeXrpKfOWyR8adNL1BnxmCt1r
g2Xl3TLqSXhRdUO9LDQLEMQDXQ5+vaRx8CEl2nsn383Wjeskmg3ahODMtZX5V7q9hpQ7Tv0gUE9q
8FdPDGmsjmGWhhxlSR+LfG6kDNsEovN7Nq4CkQIAQ2RAvddnh7CbJ/P1Hg1ClGWO4FrVF7WqOZbu
+oo5JETI3USouiiQoucyHPQdEoc2amkno/JsJgRpWEDDEol7Q2iRYfM1aLVSOrcrz+uBWGOWPN4t
it+B0UsZoTk7mXf4KNVggS2zm+UbtkHjW4Pfy+pKOZbbC5PzuaLAaL1i2Qm0gt8epnt68DqMVVtS
FNM0W7XoUky57XMmyzt9P5Xjo4Sje/2vk6N1LMaFblCAODThKndTLdxLg2JKcNKUv4Js251VQ4Pv
uKocyijGRlMB2TfRSsjhe55qVI9T0M+ToEF/YItp6NJiqk7eEjVYpBwDBpKJmpUw8vZcA5aaMn4b
08qBvkAX1kJHwmKfPzjmlCsgbi1ID7yB/GnhyDpUnnUPrYYMyizMgckKB8EE8QeM8YvdUCPciSsY
y61LqTpPniTCi2PPf2f7rYKXdzkj/ufWWWOnXSkycxbURcbQtANnK3VOZgiht4/b+34z9uC99vsW
2GbwsxhCb8F4kuRFgf6Y5NGOQd+Sk/OYzXicLjmA4XHw+958u3pukNVH8lDYX4Mq1XsZQPiEz6MR
Itv+chnU7JkeIKJNdRwBx1AZyNgmDT+ZVRGasocOEAfsevGxIH00uTiwrTiEkz9CqswIXyrxS8Tr
zhZ1PKhUWPGTa1QlIX5EpwEb3e8pm09OPT54QhYxpAfV0SgKWOSzG3t7Zfg02Whzfe92yHzJePT9
09cl2AAmVYfO83IVzQoR8O/Y8CwAt3H2X9T+5MOF10TpKLCt/Cm85IZ2DW30O3LrXH+03G3cpout
wUjkYTsmNtb5y7JSsohVeFG+2K6dg3flfwVMu077dywWifFwtYhzamCjdKqXsFWQw1R7ShYKpohk
HlGEWtEIC05BKWyKXyaI2z2D5jDd2DpuAGQt7+9epsHGnnVezmUFPA9CbF/+8pP72ItqV+eCVIRf
vJdYw4s+xZxlqpSXfYmGgSzkgq3JPdbUp3+kM+vX+lDg3Olc1w2A57baXkbamLhhuUPugkve33QN
63ckzrzkZiHQHC6wioBozRwucleF5SldQ0Gk7YSXMm7tAQPBNGtk5r90eCQTIV+r6fofUKayim9H
k1eTBiPuxy1rOKapeY/MCo8Gy1ZadX2j3HwmKF+4tLmR+cxc4+3HmAhgjL6Y56Azse0Tg3PduyR3
ny8WU/9lt5axPgJpawt0odPw5gELrQJCZJMvFtQFrLzsinjbjOLuVeYs87aEa9zn+pTWKNHblCZN
BgIjJacbCIhxySmKD73Iv7JqOSfcfroxhCNUGv1mYhgyBQOMLpptK+wL6W4qI/DB9W6BSX5EjeDr
KKlJ79OwBtUY3jPalVN9xNBh2cbAqGrt24ak4C6uv2OFY+RjQjw3tTYuYEy0K1yb+C13Tmd2nlUI
I7DTjZy04OgKgBnub6648DG+l8WNshQQP1KNcj446os586EwgKaTt8cgnkzWwnFsu3RZWax5wbCi
f8YMReXAit8THhCUK9Pc1n36Evdmp53TSksKpc090eWmuxf3zR7cqYxRE0ISUKfAf1kGWGjiNqaJ
VAi2oZSbeId9WYUsAl4UuQNy1QyVgwwl3j2WwrTsSNvTCfvfyeyjxbdpZT2YscC6SRrt93+kupqS
1s5qokuMWRldFUvg2JC5opqit0jQn0Pv9PW83UmaoWeJNBC0x04yUebnl0Stdk+9+hryhfFOLj9b
v9by948lCJEH7iYpUjnsAlGoLdFSu75xaQH3StONMvzkvbvPnloxu6YUilkBCy1JDA5dg1CcEsVN
2hKAd5v5ncLgV2dFBLPPixXtscYfUyqh5qP4xvBeUTK+a/a+Qg8v2DNxt9ZMTuGQDMayLC0oOGr7
GeJ6mUzQz+Yo9i58nWG5SG9+5+U321q4zDHZUdeuDDdMT4xk4tVK2dFWo9AzwPOfbS/qk9uxVtxS
KL1n/LhFw+x66csNoE5gJgmAS6uugnmEzFrmOB9/75BMqQZW2G4mewTqrQmqpC6pGLXNx5qT3MK6
F201/xIJzfrS2XMLN1jn/y4Xi2orvEBMNW817oY/+haur9KIEUvJUcSzlGLvOdpAhzjvAXadtSgY
i7sgsXx4F33stb4Siy/bdcB723GLFkAk4D5Sf1AVAxoPtCFXAxtIGk4BTDNVuzGBR4+bRpEzZv9t
yNuILTK8qW+NzZE1piaEmoB9Gpzl/8VayXb3ELd7zN+8ToG7kb36D4uDJqZcAQSpmiNvWu6ti8W9
VvFnKAd1PH+5SudNyRwJn83Apq+Ux1P1Q2XenWIq3qeCwQ2q/2t8rrMUdvtHwkRokgrVhQbTAqZm
tvQv0nOf5rR2gYqwwyh2kmcNS2jUWEVmR7qVefV2X2a0FGEUf1H5b4aLlJBn+5I0lPDERPHxSBPv
N/QHS7vwqQ9hAqzxlEEKxJvs45adHRhHIOH+3D9ZspFCM6701EOQLXB3GPHD2vgoyGxXvfCBfQIb
x35pbFFzcjyc37lTr4RpfeSbED6Y6fVeQ8jbYfswFpjQ/4x515B9ITtVNgQR02XGwHll8Jm29fOh
bmgQ29xPhdeXIdkWS2eWrBw5MqkVv+eTeEy60Q0WvrKPCbgElheVutQP9rbRn0m5/CT6vCzS6ib7
3VBsVDR4WaKtB3yTZfP05IRKfPJLD1ZViQ7hitDnKZhBnMS59wnk7JpMZoKO08i+P0LKkypwh5ZM
gRwWjpV1RJHpuw2X9eYIwUoet/Y/MGN3FTVE7IpOuELclQ8QV5W/1NI1jxtzh5T8KK4byRFKeo7P
A8+zuVVRE3FjzGhhBSe/98H3egiw43qjedWc90j+exfnwm37cqBbF18xN7c3rwPA2+R42UGhhdu8
kAzIi3UtxJ1cpjO+VF2MqV+kZpJgls9f7gJxJRbRxldWQ8A/SQFYYKflzJq+Fc8YycbpARdkMDh3
3KuyH1Vhk85Iwyu2/GKGsC78+YLuPvXdendhK24V9yKyVaIsr3LwbwRixzGrKeKMZd7QeYUf3/e0
btcLczgaOeftMOeuMwLpJzZeUSCf8MeNcyJwoYtC0/6yR/N5ApDa68zCB1EgLpS8WLEZoDtLHUvs
7NsSWjx+gb4cV2J+QlrnEIQKmn06u7QAumikH6MiOtPpU+VUHtjDKvKIC7pKhlzLL7iSbi3uSabU
u5PFuKhFGcHiuW+21NAEohspPteW3aTyygGtl69E3d+AqZP7jvVlCHZaItL5imXoTLYuB0XaBWO0
Wsm8JwH5+dJYe1L5WJPmfZZ7ptGn5vujxnWfn6D9CjTD0hwcSa9B4B62ZlGZuD+lSV27q7Ln4DsD
NBfj4WqkjBWG1Et2mxFL6dK++CfiXKqwSpEyziSlydXf/QBoJZebUiYMjdLMyRsHGIojTRdf4vA8
QTSnu8ZYLQ+n3uv2Lkp4IKoDLfXvnHgMAn5XT7gDvWUN4u1nZ5PJjhy7Uv40pncm3L+ot7m8YcX6
VI4JhDFkHUiHgt8XBpXDLCopCQZy1Ijj3lKM+CNK/WNeNxrOgkk+zKhLH4qNUQOsFplBMLgGPzro
6p/VpiTpeeTwyPoIaVrrHY4MBuHDYZ2fNSbPs2YXmIDX5y1J4f+wsUJKhMAmEiHj+Py5xCu2CVCf
NVq75hVunvzf7c2V8I2SitWJrMvcmzuzU7zdam/L4TDIVzh+2YwsdsVDEuE4JDD94emSp3p/JmWF
0HhtBUOpmVdS2yeF6Gq3Qz1OWRQwe71bdPaDxFkEStcSCjKP1Ln/oJGYqzbds+FzkPXG+36rKguJ
1+jFcvcY2CeRCGIgKRHyk92b3bnjCySya97eqdK2KJbm5YjmbSvYbz/ERb6e96tMdLLIA1kwxGbk
5Y1PVPIg4QMYE3GuH5fj8DQbwcjHMQEO8Ish/2xkpeplJv7JPRCdDlHlBS+cwwe6BFDwfK92Ot4w
bTN+xyenkJKk38AwgHViS1123qXQu6kGYSBwfFY2wnXl3xtUo0KF7zV741LYUX+RNnP4FTjpXgcp
wpp7WQ1pJoxcIrzd2J0hZxdDYIQ5fGv7vo9p1nHimOouCqvM4OuVtGocNGmr4c7l5cNmHRKGOKVx
zSZnw5nCLbBtvdqnDcyH7UoC3vrjY4SO9g6iBNLBK7VP+yRC/syD6cv5plUTC/WNaI2wp3sdlMGI
8cqV7L/twBVr9zuTq66hD2S0u3C4bs299hfzpIuVHRV5kOFCqXoT8h63kD1IUps7jPSG1/yO+4B7
556uAOujcNtIP2vy6ripvjSGKESNgI/66ierGXT1df2/AfA+s+QzI65HLBKrvAUeGTKsUI++DahI
4h89ThFAaJYamCEfD4pJM4Xiqz8vCPWj//znZoa9Th1pDZE5J7C8i3DxGhLD1oIquyvDC2IKQYyH
aU8JJ1MYnAxP3wSBdhpvQ1XiEnkSnp4g1vh1/K8kgPkCulmHUF2lRfKr/viAkynCqQD/4T9phGoq
2j7y+rJY0ep+Yx5qVw26aGFoeAn7ZDyFXdUYKB9tMGCAzUDwfscKqMokeYv0UB3XH84RqaX+oumZ
MMPGQb86uf87AS4DCoKeONa5nhxAFIT3dxY3Z6H+jOxOsNfAA8Vov6dIjjnqE4a/Dn31ONEXPQuo
2D2sll8DN4O3xIyEp+1c/uHHGeYVnEUAzPiD7op25Gx+c+yJkLqimGyHjqf5LPdq5gSt2g6BlXUh
CPyHnovt5UNAlNVijbH2tkKsovgC8kRjAVNpYx+M5rVGu6CnKHydSWS/ae81+wYExNpiiCNedrzn
v+5HwTUEL6wGNyTiZNrPOcyhCkpH0DXbE57ODq4He5GnBuHLFJVAi5//+43Ynnddx+Wn5ytvjogX
xvMO1oh4xshaYtWK/uX4YZ6O+u40Ht4IFRHBvWDOjvST+Mc5zfnT4wU+w852LkjwjR7rJAHkNf0B
81DADmQ9tuem6fs4vj38KbGCGDHSdJNEM4eE8eB8nlc8AXDO9j4HUDntkLX6m+uX98EyvAvJFsxf
fQh3jCM+NbFZLvbpCJf8dAbhQmhlY6G6JQqQbNfs2S/Quz2xys8cx3gvZ9gnGItfyHAoo8wifuba
YH7DrXUNv/BCEzpdCihMViXrCD/6zT7qOusmh8ZLnFSFYAune7tM6ZHEfgO9JY9XpxwhvZSlI8qJ
pQpfi27ZgJUuf/+TNjGG3CzOCgR3PK3BkE1iFXqdfP3CvnkIwM3lZDt4UMXUFVWRoG9jlBXM4zih
SPf2mYU+DNPcR80dAaAT8g9A9YBLTGgiB3GV87pG03PE7IMyfd5++pi/IJxap+9nfit2JrtWJXLO
DVIpKJlDLe//tioln6XElrfnP9hScaQY5zNqVvz9KNHuyCEjYif28cHXKqLAt22Fmf9/r0LkxdPa
nJ1Ob5DfpmSXLzjwSJ5jw/AKP9SaIQ02eAoF20BIvAoxoAt8jGpzZbUjaSEpkUOcKZ9lwHKC97pb
dkow/ukq+WF2wD69ZGb7vwEx5DudYAwsPiAfk6j+oAa6dw4UMs+V0yjyh7BgMBjnDaQD10tP0MrN
f7pkbMmO5H4KPLP6PMRwLbxSfxnirdkHWEMSd+42cK424N8VXbTU7s68I0xsPPPG9qwkt8pQ2wCE
GGt3/gHh1Q4q4Ahw0oNREYGpm+ffn0DutngvCXAPA16iA/b9CiXN1EWGziH0iPqKNcgmZr1txsyB
8MwebHriD/W+z/2Ko8qLGGsyrryl07eJUigSsldJE+1Egpt74Psu4GaASFUjAbVFbQjJNybEDQ+K
BNnxgetNixMrASckbw9TLFo3gP9ENHXWBiep3ArTO4OFjKVlxcDPXjIXSEal7d4zmykVbML9hq2w
1+6QxOqiOk4DPQkrQ2JrHYMbUvdW3QsBg9FCCLUl3mIRgWq8/KFZH/yawAoTzMFyJDvRBLHA1MTV
dYwc+jo8MHRofnJV1Xjap3I5Jn8X8I/jXZanMGLE28nw/oYqf1nMTsdS5zjU66JFp3Cm99Rc37Jv
Jrr7ePlrsuzU5alutp17J54/ebFFieqId6q6ZGy8M3NbvQ2GrtVoNYIluCZjjNWGRYeuQqw8zoJo
PmRiThaDo9tVYWhuqMIQKhi1Ov+rmuxXeVWpdAHkxDsHB5M0S73cYuKq1jYARE2tgPMyFOAcYNi7
QVXoR0ac8QJU37+BwaUN0GtKQBDn+42sa0ck4wA31mj2qo2GQ7MxHPdoNXR8TCTa+6DCUvhohKQ8
O9hOCP3v6Z19t7Xm5BNwxEFEcyj6aKC8EgPozqFv3BiVqBUup7i7oiGqFOReoY2KkinEPrm7gyyD
7L1tANp7FvxXPHqWNV2PwBNKzMWVvUF57RXahQyrbBy2VVJgRkT5QP3yMOuzEg9JJxaoNwl3Q8K7
N7+40l22mgSkLh1hYn1P5l0eVZwMppYVS3cCX9zSKX0qgoDZdv6WFJ3bDNgWx6dQRkw31roSNvVh
R5GNn7y0+eEH8PEVyQJ6oYR4AHDEOXHnWm4psYQn7kA+R6/Cg1yYa+1zzO5R8V74tp0RvxQ0UrxH
Klt6ZDFx8mFHN65memwGMeyFFNpJmBW6PTKCL24lySr1I+tD+/Bbgzrl+nEG1iDK0ZEMxr6dYLnI
2xLHZ5C/2/MbxvJnovv2ye9DBsY29yNm7uKYJDgNqXNcKe3mpd6FpjSllYPBdxFGT9wuqoWyfyGp
aLInQLoK8Q3Ov1R1dSAuSmgIhGf02BHVbCR30s7tVDkPfXoJYEoM+9gLXBiMTZQWw30/8TBpAST8
Jv5CJRQE1VSiqk0spqK20SQC1CLWwfXHimyqh6eMbYxIgxbXs4Hnq4m17pALKq6RMEWeEJqeyvhX
HwcQ2TEkqgQGfJTnvopztzPNPE7tPzmu/lYNYSqJeVX50phh/jQa6SZbzdkdzc4WA5Q8AKgSldpv
u/UaHVg9X49pyMCEPqBUdpIL0qJl+Ui5o3GjLcrvPzuGGNUrOIAfkP2ItxyIgzWdtW2ehENt6L9n
gQ2z+aPb37SvdobzTHLk/msda6TO+jm2f1B2Ng/xc0GQnIchdJ2P7oZs/ei6glQEeoWztZEOc0sl
2j/GjKnp4kqVQNy1BAAcOMUqhyQ1VRnK3o/24i1izDMh6Gtjr6h7sOsSnCvV9f6/PAUCoQvV3hBA
na5VNTJKJ/LH0TlrfoXZbWHS5cjytL5uNRbVlDhPyB2y/3+sL1Kl8cWpjSG5HjJfpDUQ4Uv/u6V4
wN58LpfDAdZmP/JtNlBPJTeCxhhLyvwM6ThyzIUnJvM17iwmeDjU65L5qYf7XtjmZAmjmLW815dk
FPGV3D4zmfioVxXpYgBeBJntauoT8KPzXmr0oJwl8wYKWfdt7Mw+LHlgQi0Ek6GFEq6pO0w4usqY
tqLA842+HLXdVL5DbpjKe428+Uy4DuUoLaQ3o/PxcoUTWNzgZaf0baSlTodEa8GGGbqzt2tkuTA5
0IRXvyyNK022r47WyEDl5ZCOXFUy69P4JhJTlz4G9U4LEIzwS8OA6HErwQw10KLJ8G3LW83vp7qI
UVB+pQYd4/1fysrX6oGjC2gs+wriEBoek0gWWhLF6xj+joPBWdsXE0J2/6TJ6zpxOq9n4Xf7t8mk
H0vGjSGuAHCqf/PNrKCJMZSgoGyc7SGtkNmV+f+j7GSarOl+GB2jW0Y8BwrshT7Yios4H+qLXxSl
5PtU/Fd9aujd9+NlIpfWBfVAdnMtxAf1LNQ8IU5DxK/z5l6UOs6UAS6h1uuS7a23paG5EGk6RmnN
LBPSg0egDZgWSJ+6B2kjOEgBbO4TskYMrQqJnFNI4sY5GIVvZa59iboCqu6tv07qjyPC5lP8pl/3
wY66YoUQDM5qfJD4+XYBDFOVSM4Rm9GYic9gRcKFldIcI5ziMcPsBP9IWRiX6i+qtSOLMjGx03Pd
3jtRqOi2OgdErptkC1pn9uToYvv8R0w6f1EUee8q8d/zJQP6ITLfQb3TrYfvimG64ehX3kd62aGZ
qAFCxPzXWMip99r6Hm6rzRB5e9yHhSGeCXZaafz0ePf0jp/rUOZVYl5P3Aw717/9yuer56he/XHC
SbPvQcR/fZhfTrU3TU7R19oWb6GJ0wClj4BaWb7e45Mg1PyLE5MZiyRapRyqZnQ37Q/svSESrlqh
z/rKS9Ys8c3sxEVdXjObGhEc+Ke0OSrQbwbdIqanCTuzDMLtXGrDcsWgaKrbivxdZNeV16uHVRlX
PlAJ7SSTA36Lk/rKUGuQ+O1V1U8HdkmE7rP8HPRm66qKcrPhhEVS4rMHver0+Bjx+2V1wP6iMFEv
R/QpIwypE1UBJKUkuDE7+yqEheeGojHy5w/4qTHy8TR+9ktvvYmFp428KTKL0jV/p0V1LC2b0C6/
Af7gRKCF6cEJ758tTDlw1bj0VvN0lv3C8Kbas310p2lAl0/+Hio903Z2QIq9XUAqvaKSk6sKR2pR
hCtWe4ipRFYQAELir41gKIJBQPMm75IZTje0nGDTyP6w2E0ePH3LyNPPnU8rdCNImf/4G/rPFoFl
q1+q8FOQDVWzXESzfsANZ1uT6o5Knkv3wHmy832uBeW9njU4E/P8cJTmgAWX2ZS2nAYfzmvXWHxY
8ikgz7DMlkrkmzE4REQNxJ1KsvrpLIc0MaAXM0gvzPqGGF+21pS0sSYvwKOwBD1FtEGSe5xIfqg3
HrAnhLVLxEhsRyu9K8CdOQq6uNzPE/KhNtu9Yiwo/z+L3cTpu4tWo4BzmrTQL/2LoXSx7byc36Hg
QhcXn+zGhHkl8K4fFWvjo52ZQXbYmR+dL+fwmRntQhf3iJKcEqCtT/WnQDYLNiMY1t5lpVKExIHJ
/yJ3vUd7sfPibL/KybG9Gi+iAOxL3nqxDmMR8Qkpk62PQMrIQ9lfUl7pAWpVnNF0q+dQq2Srqmx8
t4LHsvzMoUdHRYm+3FIiHb6NDdJLMaFGTp/F5HGtXLd38jGD+mFbBD68Af/GnwWHnkWwvqDtds4J
ntT2J6+0ptNL5P7KIFlF6Bcttn0a0ZttcBJcjaPMi19yPEYWumXaObPefwldpcYOkM1/yLt55MME
G7vDc9bSQiflwO97fDpQNr0KE/RLgy0AsVcPDgoLxk+gy2rHqKJGVBeeb03FvtSGotgZLpuNnRHg
c1H6/35jCSlapHq3gkxOap/L0d9yNgCUgbxrDZoyKYL4Ux/Hf8cuAFQS4E/o9KX4w0ec56U2CaMg
5CuJZo9S896oLjMBU6LpEopFX9dcAf4yH4XA4422ZAJEm3b1kHsxm16sN4d7rE1hFBrVgypxHFd2
5h+anlP15oq24Rn1US5AH0jiUV9/5ZwaWLj8VguZeWTAUckGi4DNPse1ZfkJKO2I4ELLjVdStLdZ
wDM7vBWn7/M2DHUHLQOVqgPLSPuDXSRgsBcr3pzGRmZ+a+jSmINru6pOtGJhdDS/pxt567prZX+M
FgPZ39DdGThCQ+tTKb0LtXUOr0bss6cvhWK1o1LOr8LT5aQ3lPIbafAvky78MnZoCOBFKcbzsNg4
dDawY3Qwty3R1L2L1wLeYAtCE7R1RY4gVMssA45fSe2hgvu8dKAG+cB6+HzrKDJRy4O307z5kcgl
HQdYIq+iPlD9pNaUb28W3MhiqOdTKlcXxX0KfkWaHchvUsAnRnfxLZZC11p74UlwpF4INIjws0sw
GTO+ULQMo0rx8cx2c5puiTkNZYMzF/Za7XpJx7s/DjOa0wk3FySj/RP2u3qzXcZHlKpr4OpL4oDI
4BIz0XyggRlLVwWwWblt5LnnFxmDTYPGDJpWLK1TIu6sSnOKcz4/u/kz1A2W86KOCA0Nn/lMnpSD
DlsOhQyxEOgezDJEd4kIn6U+X0uWg1w4SPEwLb7UZAmuQYx8k6uCZrsfRbD9D57CLzMJHnctn3mW
+BqIY3ewzR3fPAZZiVjZ2Wu5EnlldF5duNP2DobdbqyTehtFsmgz7RalaoLsLuY0ENmBm+ySDM95
ZIFAGatuw9tGOrvsEnB8dAXGWGZuixtakJtSOQIswHW0Rne9kR2hZD0DUTMXV95uHevSFmZqfV+S
2zskRdK8T67ave0B0sf8yZSI1CE/bnL30sMqlBLNe5LY6+87KgwWxdj3xlhacEt6bBnvcxaV5b8r
u+iA+W9Pn7xLGGQZsTq3xf6kqNbF3geJN4M3MfxSzQfoHR5ym9diTF6B2cjBcps5bF5BjpFpK0vD
fjQ1WayWnwblZh4Yq4Y/Zy4PYRO4XJ6Mb9dz/7VfW2VJQs3LSxixTFdxX2vgrR1h+FoFy1GLzIJ0
cxeZHLHBYmCM2hBcGdI3GmURdjy5+qxsN9A02k/4Z7zx3hTDlR6CZWSOHYDVpIsFSK1kpf60qntp
w5ye0pasRfoS7nQGqFW/RMVpLbkStcxcseOdNJFvRd9s5bAhqePxPmOfyqDY7TJKnzmU88Zro4uJ
/mxXUYAoCkUo3cGel5bVJPQM3mceY3FwXdv96RkVMYc8HFAIvE25bAAaSG3pOyDHoA7bmfKbt49u
xouBWYOPFu/zLO0TMpeRj90J5lcN3Pvxy8/pyBBPX799DQbl1QBhjGeYX7mDa6d5ZIUjnKX9u+XY
6V5aLtI2V8WhFHMqKLD5aBB/Tr+dIPWlZSoMLVk+8J32qLXi4zuBg1wtQ/IhRRcUjzmgiuZfb/OE
Zn+Y/kNoP6+rml14So/FrEHORgCKhI6RkK44gzbmRYpWkjkEs6BwOEbdCOUYw8SAZQF9FPL8u3SO
zpNsxurx87C1k/E/PdJEnTUJZg/pqhPZlI9yU0bjidttrUGcbHcFeb1sBKoNaIt2zuuC0sC7NBxx
xEVRAxI7VLQi9iVT1ELp5ikSuK1vG43J/TA3ZcPnVgeWWtMoBgQaRmoOIPuUGaWjh+ETAm1RnpDh
KS9iNK7bLvKdb4HrRqd+IprPMKQYnzSILn4gpSvzeRpYeBO8tTVZn1A7IT6PniRMmeNDOHX8Nfth
8mSBbkTMskU+Z26vtiBUxZalPh4ZOTTisE3hovjSwgUu6t6I77vJCMFk93ghSaK2FEUWgDZRb3YR
0na/1kwmg/gC/UB1/EZSbg57/3zS05gWbNUvxRjOWsmsRzwuHycd6TC2LWC4NJ9oPqJma9hTxeqw
q+QJU8jMGMLIOms0Xjg1eiPhv4HncciGPXYvQsKHWGSWc+A8rl1/VbVxK4piVAEwTiGWPwm0vy4K
kn2Ps4kAD52roQ0uWRaV61mJyffbQtfDixVoJRtQqbr0P9LjUjHRGST7D2zz2a5DhJf8bX/WoXxp
rGDhlIUbBFiJhKoU+HGoyMPQwGCZunsPYSLRok9+RcE5GDVwc7aM5og97Fov/XUPJiuR36IiOC0B
Ucset+kwLauWe0oSQ+d7bAKuNxiw+Jq0HA2cMfPIic6Crb7owizXIOtK3VM+p7a2k7R05D1GvVkb
//Fjj/rYsLG0BpJYMCGFR3J+kpryREr1CwPu8qeXDmjbmBfhP57fgs9wC7Te72Fx+TW7Pd7kt+lK
QXBsXiIghLV9L0U+zNzEHNPlzssOZq/q39v+xyddrK+E+ZWItjl+aKUzypPoX04KFi/J0Qp9hwq8
pSdu6PYrHMMs1mh1ImFyPd0AK42wBIFyRCXFwqgUTJNfx3waT91HTuZYAu8s1/rA6+tNc1lSktX3
0NAYyh7KwqHEVjzixrRNMIWm9jGGKZTrEakh9Lnq5QFCQEtfubRKVK+lHsOtmrNLP5dPlX28/tnf
+rzlGm4ild8fELAtZdo2cPGa6QsMO4Mr5BfBAPNaC093WMPdtJ21+0UiUMfnz6993OMUhvnicDxJ
Ls+QdZTItWvIH7V8ql3WCesSitfTw/0yY4VXeBzl2McEgtQQm9C8fXeBN8sWU9JCrXDTfn8lrJgr
7w8XQoO5yoUqmA819YFEHsAR3sGjliya8dh87H/CFZBZiaPWJtQH9T5SO5gnZABH9sjT3O0TMnnG
6+oQv9op2BRcmK3RqtGhPiwbW210HJ7Yelh6gSdSjC/+NfG0C3tPS7Ej7DmKqFV/PltoUpxG0Y/V
HBG1S3o82EZ5PZEdiFyoG74wRZdV9PGTKRJ8JjVFml68nl9A4zyNHpmKiTu53ZUotoBbC9MQfsS9
shLSYndnt551r1zUwWwymDuLCbTpMfceMOATudqsrxcpg6u4vf5XsAKjOM35QW2IAsM9TRIECrEt
wBhmlO2Uam/DCVGsN7s77JJBn4m4zgYLtlT86Q1LN+IygpaCbaRYuo6jOIPj4pPHq0ri1VoZh/Za
XaW02e8O+BdATncGCZsFjQEtv53jqIXTVGDPBFQC/822SqsaUrAoJQLUpggAFs761jek8wWkvis8
odk4uvW936xGOT5wE4wDV3BY5GphdAXTX9uj0jxUZ6meRDUleXF2Er28ZT0ZbAHMSZJq/RsZhEw0
yPOaX0WAwXJbygYFzNYSlAZjZ+tBew8UcBNo6L4ToUF8UKNRz4GCV00n8cdxjkRmh0Vw/ZXy4DRp
TuDHW8syYuWxaboRxkscaVFaByLQbDAaKnGxJiEzLtDKtVAzN6d390E3yedw9DXQuc0SW2YTzm1m
rKcFQz2ZNMjyBN5m9CpSzFK1wOHtcP4o45AOfC3UOjv+IEvwhyj1gRFz1NYPpG3QDwmgWdJZ5FEf
a9f8r7cBSAJlF5DPHMtveyjL1zmf9XLxxh0yreYQswn7C6e6JryekCy+pQnwkEnlW4vTw6YUa3Xv
4W1yaOCj5M7aktkAJMyVX57G8Frtp3pcthfBUypN0ivwttViW78WKplhGoRlU3W+N4dlHu3S3wT0
W2OsIYwyMyX1tCq+18uzUdyK8M5v45KZO/eIOyZRzS2131BSZ9cL/m/g0alfGR6DNbK/LpcB6VSu
FTtD+hZhhrA9lh6lPHXjrJFKrkuR4zaQDe6HxFG7e+lKUBz7Wic7dR/S2IfSmEuGHbgToh8lgMnV
nScHmrDu7f8MhSCSskncBR3l7h9/OojYlr0PT+AmzQMlCESAdH632hKa84NG4HK3z7E6VVl8X+Aa
8qrI7YgJxdtu1kdyqww064224SvwA4Sppb0qkUel/gFukM7k9tYpSxLBf9LONF4PdSf7nT7Dmhqr
rD4xuGDsplGCvhtt6+inYbPwPrtwzjKfZlJVJMEysiVJsPCrd7cxQr9RpHPsfT8ty9a4peYfLSon
iO6nTO07nNFApr9tKzlcEYWysmcbTgNyxWiX8ptbe1D/kh1VmQCaQ+ixIYRZj0wngaIIsYqaHc+Q
Gc2fb4GxU3GE+2OtdKHLJcEq9n/pBA27AmUC9vpE7xJcu8TBDBdiQI0DjVTgeDycbcVAzulYHMQ1
IDKZAysYePu72BHamP30OKqK3NflLDPI21RcMTypcgsXxAyt6JrhERfo+wxbcFNJ1/ECHH2+f0Z/
hpoG6iR1E5w1Dou8tOCsdhqxCiC4yD9N0I7YNRaSIjJL7JnztHjK+jobMMZJe5aPYoDCh02c4GR1
CJ4dW4BihNGSQGxB+nuxG8rkxJ7hETrsHXQb1/VoBTTmRLjTGysz/Z9msfuKJlIWlhiSDtCn6fEO
flrk263j0PVGoL1c9GRC0tk715ybn2hNqQWBu9Zyr/rMR0vT9ZnOcr0Pni//DhmkkiXbVYqTFKmK
ZkCsDswjpYElaP+d1rf9fygUKf7Vdk8XHHNPlZkAfOPs6JUWbuI3cbDNkYg9ZFaabF4xNeqE0Qd3
qDsrTTbwK4BzR73haVFmRe51OeUkclN5ySmJjN7IQfV9icMFvv5waoNlLb7aaOxY+oRvB2eaVPMD
Nd0m1eVokr3TXIcC8v4gxM2sFcoBYt3sjROvUMi5/s8sRE0tHtEWMSzSG7fytGYmxn/oyB0mXTOC
g8qV7GGdl8tqKeB/Azu8w1ePTz6nQRcF1fJuczVZ7l4voKdRAo+r9Fz4tOWyxmQOIUZe4iciPJgt
KVm4l2oXuYadqvzB+9tgFr2ADjWlBgkLTicNFYcPl1WYh+9MkD0Psr5dkqNmV53IZQg/JhXfWEjx
zFICDzerIRBRTbltylHZX/Op/KiLkKDJcqCBLrZoXkLzVn/f7uFogXCYx2JLaeJdrzOzh4sdIN91
E6lT9jix1YIjFVBs9A/Y3cfZq4qFUR8lDJyuW73C9FckiZiLe2x7Yy7B8QzT+Nqyc61h7Z4G1dr3
pmuBYyO6AsuRpbiK3q8NoLAm7bEwrPWfAwmP3n669dPnBQB5ojvpsDEEJ2gEQLt08QVfKLty6arl
e1EQe4+KxXnfi2lLQ3aMWffTTxgS3uaP+7eLAt6JOD3AxDX5e2035V+DvjZjgv8RncMXrTcy3HJL
mabv4YgJFOAOT0ApVEAkN7wVicHuhLKdrp0dK1REvTsEyqdiQI3tcFfNpyr7iKccXW9/nr9wmmQA
PxqCMXyYJHGLacQGfWiyedxInTVxVFKTfPSxPK0v5uejWqeO9IEuQtNDA91loT19wk8NVnXqQ3cq
C1ftuiIivVzoEHG9+8sJanHDLT3Zz4KvQksVo2buErQbiQRltCVFVT3+QGcqkPZnP8789CBe7Y14
oQg/p/OW1/Ur3rZVq7bzh07B0W9m3iIdL1zZUuarXZT9ftt38pmF84XY5npoIQFwoRAwcN2lgdUG
DG/M0OpaLGVS5HgUWSDGkEttBFx/JacQ9orL/9bCQZgcM0InFi9xWAUhxiFzu1EAqGOvsJr2juMf
wH3UBDZ2/nnSCeVg846b/iQ1nhFC4TL5LgLsQKVZ/yVVNqkGhjJ2CZPxz7mn1uQtaYhgOZxtHlYA
vZ3Rr3kO7DmGnR7AsHrnnAhS+Z8PZ1pC29M5p0EjLh6F8EIaZSQpt+c7yYYSqXCmenulTXn5qExZ
ehZeKBMRweSTvX3JoXbuU6o9pmInmN3kUES1klT5x89Ko8vCylk7YvKKIh1zefbbai29i8DwtPKp
UMevoq9tRhhtaqAFvwVrkMQluR+96TbOVEl8UiMd/vRokgScOyNozuYTxv+MdbrlCTGl/VIil86w
Fl5VfBeAm5icp+Enlbkb4l0i3P1wh04O4p2Q6eOOqYDQAfzb8WB3ELn2RBOFlYoTozvkYkj/K+UL
g5WgBZeJehNq3MQEzuEjxO+095Rq5qwbFOU4cMCIBxjDYWSYBji7HOEBs+RwgqkcOPZGjDAaInSB
T+geb14bf4fa6YgjaYJdxrnel0ypn73f/YxOQ81doeMQPx1Hr4p25g6QKjj003+49jrTWCg8ObGG
ddPwf0CYBH+CAgUTLIgkM8eCV0k0jIMqQmrDd9yDGc2acWDt2Y33kP2FIKYYp3gDtEIbPdW3+3q+
SRHg3vBzohjIA2Dn+2r3odlIr67aSaJ04NmD4ykpaEHfHyfQ9TBomwQoiFaVE6o7BRoWq84RyU+7
jvVVRYiIwH+qj9D4eonUkZdpwATykmBEl561jV9xmEEJF9+Ht+5VCcUx36cCHQITeLKa2oi6yxS4
5QRg+jPAEG9P6HgJgZvBfDZ0Bb1CiREwbS9UNYlhzi4oCqRKTjR9hfxVAQtYdoSqLpJyV9459vZj
BrYKf1jYcraJygnBNNq14EfJjceuE/4Jyk3rDZZfsNDSeKF3B8qyt1NuXFoH1e3bH+cGj6DlR1Ju
UoQrqOeFATYgu0vJU12lQfDZ/AzQIWozwKVGIn30AVLBNfF1eD7ae5kCXEr+UXapcKqtqpeAGIes
2l9B2GEyM6a001rIpEnp9zIGu7bjOb0yy38sDBHEOjCDKmIqy1I3m3be/mDr4graRnSI6DVcSdU/
XpKeVlO4SagvE6WhdzdFOgoScatTKj4nmSSIjdNENGqfnavkIu+oIHnaOe7Ev6F0LpEAc/RqZ4UZ
MYvwNxeXWy+Lu4lX4gYGZSgvrHMfvnqDRUeZhJDKCgcwIn99+at39P16O4+o3tvpuElWlBQs9laL
tspTHLc0fP8BMzb+gc670iRlXCFnP+N9W+IJJkELp1UdEQwdGw8pr2mFmEQ3hq9tEXN/jSjHgdPt
vOjilzoqdCEcNCk7+jFijM9hIklcY4x8twWI2j/AcoYSC3tE43jSQ88FrDvcCut5WArSMN9w4+8p
jWEWsovW+hbEORL1HG9xkNahBQFrAdCLNTPvKX2JqAm37UA+V2NFGXEOzGaAyfuRdAYNOBK8NoUW
+dQq2dVxRk7SaMSpOqN8Ye+M+KyBObHJ3qXfjW3BzlAmiGlpo4/o1BvLrgS/NxeN6b0fQZn8aDKD
vyRN9m7kWOX3ko+Yzilah9+cpPj7wupYdJJGJufkZNT1NN1E/evHrUTCvNew8g6PXHR9Zy1GZvmy
lGn0IUvP0P+A8GWUkA/vFELv7xjRfXNz46gNaYpoJfgV4HcMdPzcsdoJscG3S/ZGY+Q5JX+Dl91T
7fahlPJZXC2b/cI3kAulHPaS8Fn1kjHMsHkPB2uTupGz6dpIzqrOy2d8k5iy2vlJZnckItvZkPAg
81x25bM81x/Zyk1KuN0pVvHUn4Q896YlKJ0qIbNhZDqhgOybpz/XuLvmEs57f9B4tqvgv32O+dNB
an5NoaWAT07q2qAG4GONIZN890XxpH6oEC2Jbz/yNK/C1HsgvHzL2YIIJPNFMBBLavuKH7LYfkOE
xJn1X3KowQ8wA/qVxfPwijU2V0nipLyKBIoUVAPmMidEEwEjJsNT5iVuGK4hu+6eJsz9RJAfepfZ
DEjgYwRYKoqiLRyomel2Co6T9xvbplBk6U1mab9slDzXwOPHSxzUwuMeIHmBMQccoby8ZNs852s3
qpUgwHfrNMrteLb0HdVgoEw/EXw2VpClETdO8V9bTHlD5SGI1bKQa1vaAJ/498LYp9KSb34VXdW/
GTVRVmekMk7cHhf+sWowyV1L84drdYmefOfQt/3hxF2+gjNE3lwfohzZLi6oMrfJ/hhnLv2i/w+f
KCwjUiIYVG+73JiNkkRq6QSaIQF5fSci2uI2KxEDyn/upP4t+Qj23bvMBSrObQ/wjcNLHZkgToIQ
2/IQm5S/GowRMKHUylZf7ViedHNvG0cuY+1UlnFoCXFfkciIuNcfan9OUFbSYgpZkZF2u9vT7qEE
DLjQPLH6BQxW4srbvZZfbmfmzblQCDhKWigFqonP4pMrICg7O5U6Bcpm52lkqqwPlgZInlNFISuv
wQd1CRc8C9ONbjTHL/j2MUDAMMQoZdDz8seAuh/9DPkFQSD9/KatBZVyDoudjjU+Jp5q/J9qVEhQ
vMGXtnI7nj4VjDUQ784ckgUaYtXwE5AkcL+rXbkB2yf3GKCH4SZeq6HCOkNKFSjpswAWEoLIh3uu
4C1Hy4UnW2jaYZGuxX3RqEu3CiFGQlENiZ4/4M1S4hVRuhesrGf1Rt3K9xHpUvVl75BBI3wSx4ii
w0dpfHGH6ZrHioZ4KXIh4VJcQBvmI4BUyZWr0LC0jA5fFKyZ2Jy7r2432N4USmq0DsCxf/LqitRY
c2ORGaGIeHGdDTZm1RXL1SbonqRKToVkx4mBrSspEWGkauz4zVpye4GNJSZs2IaMZX9LvA6OE1ZQ
MjRhHDLSYHnJbVfS6m6X2gnkQKMYQZ+y/2kbM8x20hKs6yCWYgZk18E0lpGteh6HNrVuAzvHy3qC
d4ecLKpsvULpAjU5Y0/r883jfKNd163Y+0DrJhjuZu3dYnAa9Gxvu6fPt5su7I5cdwt4OSDahleU
gyW82E2q6YL2gKr2mLcckREWdmZ4Gt2bTIdBMq3fnVgHlP2yJbEAmh3y7saTAUx5qjtBAExfNFIG
Ji94LZ+AbW4y76Oe3r60OwuU6t3OkGlNGgHV4z1vLt/Rhbh0fFrhaOLD71gEFtQPbcbaR8evZji5
ci7khIVC4i+UZRR3/+UrcImPTkgQiyJTCpR/WN59+fcG/WroOynDvqtwJvrg6VBLf4smJYcYvwMe
nz3rULdEajCxf/AJHwO/DOqL0wcC8N/2HAnku3QP7aBNaE/E0XOl6CN339d4Vql3hXpYOyZ6genW
digKF1lWBd0uUAfl0piH1ZQJk1GZxF1RRy6mDjklrq+xRQtvqeTMygjoJXEfdaOYjOwjwDg/wLeR
qSpeHOnljPpvUHgNANrpiALI8rDqRZO6ODKTjh+iPE904Ex9GqQzTYRf1rkEVR6BEtC90oqZCMVr
1+vEzMEvnLr6o2KS7mVscRSOnPRbE8tmZ5bm7ePPee5ppUciar/hZiDQuRV+iYBBwY+EoYEZU9vj
x0BO7n7fRPiIbw1UJoPth9xxA7aYvN5CXzDB0OKfd3W4C99poX0GmqpjEDuWndfxR+3sLb3qvz9P
/NWzRyHMNtlvCDzYmpbfYVn6mWobcalmOii9nAmm4kVXz+DHjTTlRScIr+V/ERJlqMO2JWByqLpQ
nul6ORZkg/EGh06Inx7PMH8TuPVI5SdDyyLvXv6Gc2Zq6LBc1WxJmrE27X+tDq71t84dBkHTk5dp
aoW8h0aPKeQOIblWtdGVeYfdwdt421WJcJD36SjYDCciGBc7WopR/LK4AuplXjFJuqAfeLHQwfaw
12BZrqIUN8EL4M8RtBuiODP7bWjAJ+q6QFsEHU1kDNaVR5X1sLVil7ASkhVeGgk65eR9navgE1ox
juv9AKuD/RoKU8vaCEY5o2i5KqDB63cuGoB+quFTpBStoWK9XI/f/kq8eIP/jldl9hZaE9MBsj9D
PQvtmCpZcSIsD2dsa+qExfreDqyn4+d8E0Y37UMqDUgAtRzIRirH6LtG4mUp+4u5npSciS0g6q3V
xJd3SpySe+BL5cQx4HH4aZzjtibsztpeFGQ8fCRDcorJtj7wyzrcMEl0ZOr4eULK4/F86ow3BESt
znqwtnbaWoTz+zTfd0PAXn7vsGlfqmJIU74pqEjOKRed593aLllVABxyIra8b97sGEWxWllA2f7q
8WL1E3G0LGRDkvNYDjk1S7QkV0fW7/NYWb0bTsLAawniBra8EaPxS/sZFae6HFiamdxUS14MOnvl
AP8/Au9jP11Yz8IaRM61z2aFI8cBc8snyAlknT8f9KORYqzMApkJqU4agXFCBkWX+OsYKWWXXxHS
h3ydnGqNFDIrYBQuc5wO5Fd2mKBxRtntbcE4YP9rPuXLr8Xfi3cHCPGv1UAFNrpIacPeHWxAIRkS
tpxaOJA03CVAjD98lliC8lOFZZgI64ULmZEmXaJAWE7FqWRfmG3mzsx59lGfItDpBq2S+8MwwWq3
xI9RgQDL6LMgGf1g26pCL3FBwEEnsR1rNwHew8WtHU3BErFO9d4uabMubklPFDzlykDURY8NJWF0
D/AshyYOviWyVzAwO0RHr4FGzn9oCyU+9YrS5mvEdrRQ4eQU79mIn4jZpKFqQ+NS+zbCDH669AAw
cG6DRKCBEWvpAK7gC+gN9MU4/ygnwttMn6vdlMIkQStSGVvPhvhiSGrp6idVzZuxsm+22NaZTkxg
haihTuRcBBYbVOhfU74Z7310PIceLTg8S9DLYN/7XBJf6Z7Fc/yejQomEu6qdfi81D7EDKU79x66
P99Ib+wZQUPVIoLBztYku6LCHQcD88J/zkKApPt8uR8L+1oRZQYezaFrC6ywssx98ZmyLOsVOLtw
rU84uKgyfEwXmMX4D1eGWlMMkCeKh7/KVRsaHV8BPNUM6O73G8ouizr/trO5PNqUAesQg+zjW6WF
UT8XtMhiOJ13+Lzb0blMTD4UCwU2utj6TaFEJeWN9MVq3NbbmBfyUSZI+pgjNSOAJdNODJ2Dl8y/
4ecvxha2fbd5QqWWpGaKqlrx9dtkpoKqgpIBbHBqT9arTFKkCQ1rC799QtBBOHbYKARVB52NJp36
q2iLVfq3VdmTGpYlClM/l3r0MilfSn7rE0o7201RsqzG9n5BtqdxV4bXHipm4Lcq5f0grUzu5Xnv
N8r1uaeCcdHaNgaCxp2jwrA+yxsiE1es4c+yacJZEewydJQBcnxd5/qogr0w05C7l4j1YaowCghC
6nQNDZunoDTfkL4LfSswa/PBipEPfgFCEUop3aKqOWzbt/VhY9Nj6/UalghvElK4SWMDjzQjORTu
bmh+++2/x5Eb144b3Rdo1JY5hsA5u0STQ27P4yf4mCW13fFB4QdLzQJbX1dpw/fTlNwnTzM2Zztk
Pv3iIxW28vALwISbXskNMHF5LGptaUDqJ1KgJOfW+mMjs6WjXM+pp091pV6tq5RAExDXxzqPHLe0
pR1dsW0U1G6oW/qkjGgMlLRj1LjkMPEedGtJDfRa3gQTQm+Lr0WZXOl/T8ZMwMIiuHpSsUj7EAoc
/E8kLb9xvlJFflGmQUwf0aBvEzalj1inXowJ0WHdwwXg6SkHE5yjwFt5POna/nYyltCjYlgtFDH/
yTsqDcUoRQKc+/oc1OzrVJy7tHXI19dzdkZqpdLPtiPGIMSUz9qpahbJvSBRePlXMqcduvzKQctZ
UAhOPRhewX507KZ7xFCYhyAPve4My/QrdziONIVl+5LJM0epKO+cOgTkN6Z6H+h3QgtYO8tc0/rD
Juy+gxD5CYJ2l2A4tIPpBE6gB2IN+GGygM85zG/D3f+M1iZDE1Bc7DLCRzO1tWVtWEGes9Z2HaI6
BkDz0ZfmLziNR9qwqcn3LgRZxeUkcVJgbRRY67nut4o7G0mJQ2doQ/T46sJ5+u26ElMDjWhTQ/li
4iHwDOwivV5t5llZBHjSOP00aEpd/LpbugEqlI19pJMaz29WDQCvvMMkMi7xSklaBz7x8w7ccO3J
5bvUlGvw98G6LlDXVOYoAgRZ6OG8+9mZGWIFdVa2hC99JKSiKiPZ7uSubBMrYEjQ0OvgRNimgUrS
34MAZkuiYFN8CDN+qBBjnbL5wi+M/N93iVISlRWJJ0jZNTjJLcPglPiBr6YT9JkjTJI1ZtbHhFLI
wH/kEaY2xMuhGzEcpkN4mLHVHqKWH14xvHSFBl78dRWE4mIn0mpzYRh9Qi+fmDX7t1VrRDOVtGeJ
NuCx7q1/EzFJFFTP2dP4Ao+xCKkdxwIoxOuSVzB6bgPKhBBqbyfMkdL8l6tmrRfXgTNdqXL8MDjM
Q59xARyUpfYKm4+eVW4Q64KzPweXxUTZqtoXo7YvOJlFuu3XITrglMulk9KkhhCWT+br4lwNMq1b
pCO1gZd2kjKpmIJ1g3p1Bt/r4RDLWccXezcDJ16UfWmxG1gG88aVJ8fi15wRkAcDJoCGhgI0Uj8h
8aozz8cJitVufHhjqCCGGY+0Z4w1lOxq0d3dTWIcNG+E3yoClsk8a7Jmn7xoThB896AtuDh3TztD
Pe6NQglPQ5QhC41285PL/sj84bYYtX0XBzuxYW3zpMLJHB/C4N4xgyzcHF9wV0C8CHc2YjSY/AzF
Q6Ivs2yU0iKZMBsbUz1NQuA2PPgCWsvNLFGtQi3RxaGLPGVt4Ty86dSYEuWOLhA3nIVwvlS18YbK
sqFG1WF6/Xtg7uzANBdUU55BSiLA+DftYOClJ/K+pcADM7TI9yNGccQrQuy1p1fOPGd4K8MwZDCR
AEx0M+UZEDnklvlCo2GptaZNRY/KkM9vAeyxmT7NqugKiBpkH9E6jul74LCV5sDXP1+JcbM74ewu
b19ZkP344ZFq2RlK1goFhhlKeHN1BT1ulrXTy5aVDxMgXxYZ22XRPv3ud41BtV5Ej/FUOP2MPHX3
GnLhOYJQBPKGehYJWWRiW0NJC5P7uHbcFJilbLVIhlAn0KIDIau4ZpaKYwXwoYnBHejJIgus9ucG
IJm0B0SzvATo7O11E9ZS/bSzVU+2AHShKwLq8iw9E6TGWGkXIlPptqoHuINFQxZoa4yCav8VDdKp
OQpfdhYlvl7M8Aj7blX9omOwKDceFCn7gv9Ak4QndwAzNUyNYSRuUMZcfMkJ5M1Bp4py+TVxEbsq
+jxP3U+MLP57JP1i0JzHjvIpI/8/yQnvKqlQFLzVdDmmr6iQlUGKZpDZmZ9uGx+li1zyY/6vHqtH
SI0XNnNKxmsCO6lySwAfvDWRheQICdIzN47b9ikFpqLSGSEWuXtqHOqWj8jzfcJVsPhvyl8g1zrv
uCDrZSfzGc/p4vJ+/2m4RxyovPLZJM8gO+C14a53I1RFen8hRmx7FV93lC7o4NxTwJctsxC2D7mA
Lsah0qxEkGNyKfAs5Hg7V3bMYp2u6fYf0WxpzjRXSkKqcIuuDZqFvxU9P7Cr5owefoPslYfMyDfL
2dab+DakgVr1oxf7oV8wx7p1/nriTwmDKvfKy772E4xrUWsIgUAA7XFMOK7LiB9nLb9nF58DZXyO
A/l4XiCXIHWgFVk5d51QHzBGCpawS/pjULDdSV3FaZRWYqrvIJXmAjIueEcm4Jz6U2gk7Ex0ZVOp
WMzAZf9kQbUMOe0jfG+vlPGPR5yOm5PrUrBdqGjaRBag2B5Sj7knVz0BX02pwbxbwtxsX7YIE3Nt
+xmei5gbXMhowcBIyvF1Whnz59mRQ6JBaIcVQIsWZJWE0UtUiH2PzHkg/imCJytiGR5sFxFWCnEw
vHcGruNA0SrmCW0NbcwrXm4AVkWf6On+jP0aR+7N3HB0oU7bQ0aajqN3CzNA3RXOZNhFurWM4YYL
eq9jD9LpQ5nXoLMtF+Toepel6euifvaCr3vSrHVM43gPnfWUB62eLD5rWsNXo5Y0DMZL1LgpV02t
y6iGbJl0h8ZkAwMvs6y+m0Nzz093ot6I3ZyzlfGq5pIRFdg3ZVLG26YR7VoxFTciuidF03zMdXiw
BIOBmsJa8pRTFIXlzqOWE5q+ytCYWY0XEcXKFC/63F2ui0ojRKW3UjGRQRvIvOPhK7WNyXoTIlJh
kTd1WMaG9WWi4VesZ8ULae7xZmDD+hdqfP8D0XE3sNzIorqzh5yfsqX+R9JnMFVnZ9WkWYRt3A0k
77tGTsD7xcPFE8piJji4xtwDwK2VMNLnWM+v4rKXunihUF3a5BYk19IhFk/9ijxSc8CPU4bn/OST
TQpVXvlgQRUSBUFKN8ZhbcAd60qspzgxQ9ijPxUG7wPXzQ+HPcdCDjFOG6hm4+uFt/689EHx2Gvp
MeFRVFC8B1Jgt0DcpbFVf0hIn0yPXqFUtXBvcj8B29Fyyi7DCF4x2pIcRFEGAlJ3hKtWnnT/wbfu
jJsPQM+cL4SSHV4Q2/hA//MOu32wBaczXZNsxJNCEQjIqW3pILxc/y6c61Ho8lBGzhXRU/7z2SIP
reQL4vNF9WgKPIhVzYLFoeYStvvR5akAM1hJ5V62kBhxr1op2KUtt/u+drszf4f59CP0RY/vWeUv
FAGdcHBJp4/t0VfoqUss33CD98DR4ST02fScpE7pdDIpI73JxHfAtYqbhj3n/aIetVIlQ69k3H68
Pz6rnl2ct1qbsIg7OMg8ztoHrkO4DQtA129/mNge4JOOlCqE8TnxwA0A11z7rlwq+F4k0CQFmx+p
YSwt8SxuFUj/XtsLsGQ7+RvbERDG2O8+5lZZjPKR5tIPo41nNc7hgpLyly3KHOpb+IvtM9wy5uXL
Sse/9p5jeafBXCcobueMbhGx75QqhYAGbrV3gvB63O6n1k3n5eEtyILyUm8Dy8xKCrugNYzU489L
9wCdi3uf6GfMVGUIeiTBGrpEyhUmStHUoUm1Si3k/G3pvr7XRHRqD5uaR+u0d5RbS4DWHj6CNHnW
W4SqsAKLV7jCqu0liynSLbG3MdsT45esTfV2v3a1OhAn1wa5uM6eLrFiVDU5rokJ3W+Ihu5jnO8/
7U7JvIvi0MLCMIfjj0XeQ0dBoMgQ5SNy3iL3tyScm7bD0w0WAc89v+NiPFu0tmHnZYrM4ifxePzk
5bkTvSxlwKIJtFqvvK3HKVBb4C59fSjsX9gvux6FDkmJwWpUtDCOpUXzX2Y575HjJaL6qxZZGeWJ
XWNNk7srAhf+bk93FoAwrpdMg/32cmdNX2Ywdp3mzPLI/7n8DaDGIwQqXZzOjZf29i4gJ+vr67M/
S9Xfp6NpRCw3RChIxbpY4i/tdxq/99n4oE/zYV82Z72hNNGemA8OAedmTA5u3C09TkKUNnACJeqA
R6+uOlpLck58zRgZfyF9zKyAMvNuhjRgFTKSMlGtIBxIdP3ITRJjMxAt8GkYmv2/lOofauUZrGvm
wpBUs4R0H/LVNcG+4Ey5wb//mm9KwSop5ndmdUUljWJ6oymnuiUc51/PVsmVaAy0c66IxzIYhOsD
mLHTS0BunA5O4FW0S1s8G1OQdInplG1uUS96sYa6vXaFJ37uPUwDu9gU8Q9Zpfw+G2MJK4OvXhRK
2cNJNVyQnl3Pa5O5gfgtw0hcaAoBDkEkKaElpmEodBH9sM4FWr6nq8qgdLn/A7n0HMKeeQzq/WsS
hpFIztuaFe9We9ot9WX1Mg9lRp0M3eGHlwi00NkrmmigrhxW0DmwMH+mXcKBaPmB+k6Rq0/5yR+N
0AurgEWs9gu4MWnA/L7yB0AZ4twF8mDwp70UUhjS59YfwZQv0hs8f5ekKfdFLA4gDgQ3A2B2JM7L
gUmoeVI11PZGOLr0nJAGYjFH2wFGUT/2mA/9xwbZZcXMfxoo9YY37oE5590TtDf+jMstfNZXyVu2
8cZCGPVTvMSefp0Tye1rrE+iZTbj/QDZNxfA5k5i9mz8VmFUkVJ3HShrSi73v0zWMB+KO+yZx1xd
zhDxdwVEANUD/A24nXjgeh+bmpS6fDSPu6zYKOisBDu54MCWdijwNjcCDSqTRP6EghvZonGAyWYz
dKvHQNm8EAHr37CLP/180gzsk/fyF5mIrk7rU2LASYElrLwJRI9ix+Wu55Svc5irsfnUZRlk+ga9
XNX/581jxN+JWhpDsyOGYN+FT7S+75BNpRexl9CiS+QXhp8IAzW2MlF3VQu+4UqIu4mdLimnQM6W
KtgaVNjxLZ92TdkBjdk7ulzasUI++0JiYVSYW0pxg5j8NRXK9jXZuhBiKCRRiAots5xJk925kX4/
ku9rD2FGmcaQguEu1619HSDLkRLhz62lXVJQ+MeX1m2KFAlkqlqWGyw6dP86oI8fPEeAM1g53XrG
K7nVwczInZi4hQRsUaksd4L6qzyyQu5nNoMJpHR9Gp6w5BgyoW4LdkUaQpusbcn32WSOOEr2KCUm
ZeTwTKXQpYPgw7Z5zJr1jQaQB9Mn2f9RCRy59XSD4WUI79vDTOdwYbJMGhPW/nbJdqcGEjMhP4DP
Puc2ucaqbyqAFJJTwjoeQ89ITt6SS/QDoKKqIxgnKsTyXyuvoG/N/Dr2eYuNlDX6o3IWk3cJoGn4
loW0lKeO94QG6fO/EZcqUfpEpc7vcJ6y1kIZfNk6tuEA84VPxJQfggoEPxyLYTMGlvPJPrciA20B
IjJTBMMdCOb5bGvxr9Us6dlslwtK3eHHLXA4Fj2hWQfCXYQFiNUUtpG0bPLt5G7DTxMUVsq2NsKY
IyHMV76aHBu2hpDUabqL+scYpHgTzmVj/WJFGcfGYXQmgB/O6F9dAoIh2RJitgb2LisscrFneqTO
jTvHGOJlhq7MWLuErIVb99ITESbo9Uj8GSuJGXWZvJK9CyTHHsCce4IAmYfEaUU3B4hTRujPU8PN
4Sqh1FNmfizFa8wlHOb3R97D0RUdxoHwkyEO94Fs6vuZHCvbF5ckQyAW6F0CbpJrHsN2gpEZO44t
ql1l1rBBisqc+npG4oR7PS0ri9BnMMhA9jifqDVriA4wi2a7IVpUYeOwCSjMwDAFP2iYNUfcsZ2I
SP2rmtKucSbZFVrZUhZjtD8dwKWI3FkUPnkHwgJLAF4lIpiW2XZp91oAdH8rOJsV9Lm0j/yoPiy4
YJo7YcDjvnNfd5dWuPRhGO4snfPcpIq9YPQwOoREKdl/njeuqLwIXizLPSoS4TtSm3vlzRjooNin
xeF+LzGf6G0LwM6ed4ix20JPIRI2QBOq4MiP4i/Cm4/w1Xq9lhzvKfqrFR6ynfe+uvF9VFpZQ1di
LR86Xju8r/DoDVONdv+b8q73zC5/TqTwLzaKF4ecEsv24CnVV7JP2Ss3XLAbvmHCj+5ro+nOuNQC
EM1IFm8EinvXsPnHvG6jnXsj3MtL0wxr4JCQJZofc2/66YOud7dV66PQpPkNlLpEi12fELbaMz2z
anAtqqgQ1tEOFtVniXDV3x4/BKWQ4nrAEzf3Tsm1FtQ6nc8Sxrw3/1E2PQ5QkGUayLYxTnndY9nN
Dxm2f0m5OlPh9T+V5jA773R1Kl8KuoJOafjgidXdBX4UMsmcpxMH7JMNreAzmyX053MQdadlptKP
3CF7TX1So7HaV9PlYHok6J3TX3kWm41s5WhwcDN39A5hw0L+sArYp5kdrVzIhQ/Pq5XA/QY7fUZR
LKinJuxQKVFf8pspUkqnf+/lAmyMoRKBaWluE5S0Pv066/LDBctXVMugiQFp6viqwI2pj4NWpm/x
lfGcKScBSAys35LWvVjFd8T9+7bml9k10wcSFsCP/m5znp38yY/YrdRB9fCYY+hu35nVARQ7Njne
J9B+Pu9ihEJKmhqTrEWXi/pFWvmL0f7JDGeZane1ftad2iAseGUZ+tsDNyiV8beTNM7LGmV3fNEm
D5T56PwObwsdkGAsSrHecRB21llTsdE8MQ2rL+j/gSWh3Use9fZb1VbmmjNL1FZW1gfk2e6GlSmD
8gUuRGbEKD2pkYDZAjHyw5cmkfU+ecIrV53koaKrM96pKQV3dnyOce35dLBad+S0E3uwiA8lPH6J
DsIVZzPF2VhjEHkw3WnKnC2jd4y9A8mk/AybSz+ZP81ayivT55XMlcxLGN3M75X4DcS4QRbTqwFk
REHOcrpgBhJaJk4AKriIHRVTroV0HRGde70cg4++yUSJZruMp9pW2A5fateTUMaJvBafkb1NahFz
262kIYQd00Hx76JUOgBOaiAnSgLC6LNX7w/6NsGPlzFgDin0+wBgpnbgxGpKOa1J6zr6FC3SpAnL
qe+45oOzonmv7WqKmGw3wKj8EiraPhjDekEPEPBwmoCRyalEsru/QKRII6M/81heruQFotCyou+6
0eYvwcbKpTw+7KOIco8/ScTTMbvI0E9tRklu3tf+wFFuPW2GFbnvSMhrm/e40DFRN2DqSME3ZEWD
xDljCgFy+UcCYnr2ll8Roy5dE3pjC3H5ClFOKQ5jwv6JeBdotETEa4msq5CUsftMzFz9s7PWrAvV
dNxKlzkc8CbZEFmRrBcRuVlB2bW9x6Lj0GeLJ3Fr/Gs+gwunxWoGT7PPf2yW2DD5I33oXLWJwIPt
IHogudDX6mPcInpeFDtGTdQq3Jkes5fPDhhnPW1eBemZv/HGrdcdUjLx5DuQyVtjkVGTVm1NXpyM
6HZFAJ4s/4EPsx8yIa2hKnEx0oGClZO2IL8xQwJRh3O38NUhpGTm+eIc0koldRwfyipElePQbBXM
B1FI5+j6hyCHVt3W3Aveo2am6aD2aDCeSdvccVFKhTSj85lenOLL83DMYZf3MF9w6v3MexWuLy52
+kWxq2li3q5bUkVd4GrPbc/Z+F8F5C25YBDno2NcoL2dGHv20gWPNd0lwGYS6VCnP50/K4OxI9WW
TTGrugXcd9tylLg6Q/JPtEmPqfcaMUCdcqsGOvwRo+VMWj9ALwwnlxMBfDlPIrKZ/imFOQnobQc+
vqcjnjByEGfQI4ymRBEThRJThvvoyVpKThyIF6VEsfeAtzhGo6m+/Z0M2/SWNlRLPv3ECKOapXpn
Cfxmw0yhfDTA/K4dMKOtD+18o0VB6MiLWMTrwHABMgPhFCih8V/mSDeFZ3gN1x5jM8N3V2GcZT/L
jI9kuNHwlVPSNkxE3760+37Sz7v7jsUxDgweXsExrWmFYmgsSHr72GPxt9jl5HV2LVO+vZwei51I
8XfMTGR8sB+U1YRhH2AH1oi0DC6M1R68zlCD0JinaQKCqJD8xa7JTQnV9fZi6yy/rXpbSLPFxKeI
QTQoPSOb5sJBzAlBlDTJTevTFFRRcV1eLghfi0xJesUgLUbRVtH6dGxawm6bO4VPAlQ1ruTJ0mS5
agUC3vCRoGRI/T2IKkzob9+7FW+0C1xmu7AdtNw8d/E80jKn9NaK2Jv3I1775t6pgNtv+LFdl8kq
cY8WWwjRhxC4D7q21Pqndh2RT2rbS3Er9rnrBvacw0xteOW1JkqO52wFI9YLop6yL0Icbf/9E/MV
+cORuBdRqa/xBcckarQTkrszsHhN9tshUIgWz+tuFIfmRX4Sd7KKSM8XvPqHgA/P+1WB1yo5WzCX
fiio6Eh+5yTuZWHY/g+BLL1KuDhQGibpXXmWNaDjJy5yT3WiYH8rFThQCRTTzfocdAajivReg+0e
K/8BxV4tsDThY+vhoYEgYe6oRQ1tuHP2Iyuv4JLLZvCnyZKsI1ZeWK8gkJuNTBZ03wj8C9n0sd7f
gFo9xGlbE792Ljq9cldGusR/EfmJ+B3430PBIpCwr7FcwG2HEvblLc9e0yG4BmZxKZtWpE1Bal67
IkvtxD7sHfORyIAsXM7MPa2FMOBJ3zf/gTLspP+/UTQjxGnuO3RYiJ7VgL08sXTDAmDMc4vaY3AX
6Z2sPk4nErTtvwKW2+Rn6PgUhkdAccnc8GY1ZFR6IEfKu9L3mkdD2ce4jhgnhpUeyDjUzJE66Ub4
0oLdZw/1/tfP6gA8UExpV8XEFHGQ6g7YBMYlUbbE8ZwAKjoOg7PpamyJmZNpIzUc0TlprPxcp/BC
+29h08j4n1p7vhefVMKUFKci3u0U5vaCpFGXR3Oe8HtyXzdXcP8VosqkNZE63Hyn1WRAvtkpeyEm
zNoBF+iIpcUTMEuxU94ZjHNu4D+HzyCeJAc2hXxi7EwzKRhZeybxLq/VKITc7DZtQLWQIswwM4fk
PdfbLONo7Hiwce2pZvTwzCYuyb3Ya55d7BB6RdXYe1DQ38cAJLUVXX48NLOHqj9/f/iJhX/vYP5J
NNJoUAQw8Ofd8kxar9d2AYLMC8w+EvtKyD91Tz8SP3CiVtnAte7BlEeGF9xOdp/LJuXjDf8SeOnc
ctiF83j3kjHBmsjGvlk7FWWPa2bvYDYg1Ivk48jfCbZ7FEnEUwqgb60tPV90G4kVRliKmxzFzTzn
7loeK16wk35UfroSRlJsxAOYfGyTpt7K4DYxnwozdmUxQm2lR0mmrDZV2LDn8UGdVsOtInofKNbO
Z8mRUBpzMVf/vQzva5Pt5CT1ohRuej9CI+5nmXOrbthJZK9pfRwIcigORFK6RJMXrkCGsCiXU00X
IGFucMuhZmXLHQEkVfJvPhZeeNKB3YpSFbFIuabNASaJvjBchNyMGttFMEqJeUe7Io+CX54AvfEE
cYmJpYslmG+055o3jghlA5ieXcOKNIAEcgOVGchjnsWML1UfOZS8qYJ0JepWt9ZhlXyf8YaRyZUu
rOYr1HKKMVfqVRBcnBwSA4P2czrUBhH7ixG9y+Sai3brdXMGMfMiUC04ECiscBYTvyM4o9qw+GYL
UOtTSxmHNYuS/yXi15BqoHy0r71QveT8AXIaPBEFmVSD61edlFQ5cj7ipwaD29VN5zB9xp8ywQ5V
S63ZaDm7cHt9NOFfzC5dHL/6dOr6g00V/OtoaF6m7Bp/iv+h7XrZO5FwXooGgRi6Rvx4q0E26oWf
3shUVY39FNo24ZuSWqxBgeA9rpeEjLGTzWHJbKk3nuLpzr+L4WTkKGhwT2A7lGNmwxL9n5gaPHGA
cBNR7QS4Fejo1c1pRt+VJecrYedHqnO20eWVs4fPVFwe4hH9bTM5NepMdB65zu1jbttwxlVTkllE
/wgiUjmSAK2PVI6jANWSfv1uxRwHPlgvXHtMZgPPQVur0VcT1SnYyOWys2ut85EpKIpp3eeuvXu6
DkIFygCh3vAaC5N7aQ+zlP1tdJ+4LSAfqMaj656FM9pAtc0RTL3/gbp6o09e4AQVtYRfCWX/kKwW
Ap5y14CeDdLeQGZNr6Mm2aelC/GE9Q2LVGhMb7nEz5C91ZfVt0x0gXfVdi3frPM4bZ9crhJWWJYa
agvcz3DkJSRWXd5KrT7K15DX4OXGAeJUm5Y4m5RhtZoRkWRKd2yJF7niuy5fTZVQ/NLAo3LwwSxM
TeKqAmL2bb0B6LT+pvq0M8ScjYzKI2M0sScNoasH993qV5eAUht2O45Gh1UF3fhEn565Hjorc1YV
oWdbFCPULPOM1Koyltl+VvTp6rsDdraoL4ng96rMqWzT/Cz+DxlxP1p1lV6CnqT7tyXXAkvYjC6v
jIsXKAsuv4BfrnjLlT+PfMLw2hB8SZJ4DeRMKGx5zKbTzV5RXCE/7Tvr4Iiv/2h8YPcWWjjtEdBN
NrR3AUzoWGQyxTBa7xNhLZI0hA0xbzX3J4ubu+DpqvGOM/KqO2ZeGjgx7Pa6rzzvS5Z+MG/U3+nW
3bSsr9ZOCW7tMgjCCXOVdvuNs/5L511SNH1kK2dvF/ZqnZE+kVDuhATsfOHTMi0uAT27nDOa6x10
ggnrNenjzDGFCoHfSAM2H9rJoBT8sV7rcmwJOJVyMFHLZgHo0OuMHMGDE+SjDrkuRGy8QX14lMGd
eEMOGLr0pwWA+/Yo6PVA4yfycLYgU+KQGKxRh+si/MezBfL1bLKkwrOXS4j/TJ4K8je/D6Jx3LUL
Em3vFvPF5vfTBCJBWhXBOugBdDs2TkKahlWsrb2nALOl65+qGyxzW7o1MPcLhBj3JQ4fGm1oIra3
JycLGhOC76mIbsAjYribKGq1Y3ZSY6Cd48lALdGazpaqN6+24Elyuytr9dcs1AH8KVA83pbv/NPh
QfQX8s+2NpAbRfYUAZN8PFgSSFiIRBdzmfPeXqC/gYBaGAb8CIR745WYz44s+bMwcvXcLMXxB7uA
/DCRxXFsm7t/5NCwkJNiVhufke3EC2xO4FoLR9SXZyOkCtw64o+D5a+7Xay2QX5WrvMO0HwWLXWj
AjZ9BDPmr58zpRSKwjJQpOtVMdfBPPP34wlIR0KJQU0MbKcN5h1JSGRdSyVBLoG4F+q6ps+cvZEL
lMOkJZl+0nPyrnCvM8KZi2etbONQxzSZEC9cfy8SJX2+wQT5SAWyHkZbJdhkjfshdZvb2Xe6sThO
tNSLYTPH+7CXhmyB8S1YNakK1k+5VbIK6JjdZQ7cOFedTfQwXetDjdCjFNe7TzDu66/MhIrBmOrx
lObJ+EU4R5ipl2kjFqIugQIZSd+XzIUue0Wkm2jlmGP8U6H03YTdYKrIc8szz+Kd7WqgY5ADChMW
ZJuduvVDPzqXi4/dpnwI2oeFKUScGzCYpeqzz1xAE1gIo5jmzPObh/pWNCw0VTYEIACLL7W0YB42
JCkEXeJ3u1Asv/6hYvwSLygIAHbhRZ2ryKFNz+R+U3jACT2bClz7cJJzbBZ/365w0NMFLZ05uWFf
NY5YcemytQOqSOaPNhfUewm2l/Q/NE6MAIx3q88IRkDyzV9Llv16ffR1PngFgubsZPrgJ1RcuTql
uYGytx5w6Jtidc3Aji9HSPAhYVkp6SEivCdgW/qgu15ybCfLW54IHXGlX/wvElugxsced1wgG79v
Ap7jl/RM5eT/leEsIg8S3+BspCOfnKGNCwDoJUuheyKIgm2lj6rDtA9oibg6ToOyDEH76V6/Ci/X
yGUDTu1Ivxrd0SkRWMiPZGw63QgM2GQZEG+rFLYYvnEO8jxb2OSOb9ZYG3xdUROhlokA2ZvvrMNP
wJDiivKheJ/x7302wUuDF9efVCVQNQY7Zx7Ok3O2GAyOGS3fJsXUnxs4jI5OWEM+IWFjd8cDIXaP
MywhFiJEV7X+rxwYy/E645RetiloYyylNyROmFRxJqX4mV7RYW/RdYPlIIaDQfi8IGyJG/8g2jBA
KrIBJIATBiF4JNinrmEzN4AudxWucJjRgsRe1+AJ3jqLTuZFFo7NcFlzJ46CiSMOfzgHuoU1sdOV
sDRhQ+BkSHUws/jyWKgoTqY08Qwyz0Bz49PMj3Li9vbOoenvzZLAu0KBfHefxpDSmvLCd0f+lbol
OiUl5/g+vpsG0fRSTJzqWZVRtcUVHctsJWNTtL/dQzl84XahfEhQBGjm91q2A0g9ejGOa9hXYQGg
p8xrAfQDZx/A9XX6qBMBcXLVxgzTnyok3pL8bNA6GUKgzJ2e33G/5KmrfoIwA7/vtvzo4RjvgmoA
gyBIsTPXup7H3PTqp9xgXWE7VEbufw6CM3IR+GC0YIP7+0zFx0ZMkPve1UW5wTtRtcGjdEabgiOn
XRbUxyPz2XDfjNay0SWXFu0Gs08jE29i2aYAWD/6DOSywq6gtmT//nFOennb3B42u5FrORzHG7Ue
+/327n6wEdCu6kfcOIsxeqkWNNLBgTqQ4L88NT6IwWOZt8a0FQ8WiQl7lWg858Go4Q+Qt1Z3R+hb
4x9tUpx+hkjBhDYDWTcaGd+ZTkYos1uKILfovnAi+HdGPR2foxZwpaEcIy1yO9Amq+6neZKs30ve
B7b8spCGGgbKXUu+a+qmhHx8ktanaF8VadVo9coJvqx39Jf8jKp5/ulO0r0798Sf2mflFRCNm2O3
2fqXILsjBttXRROpgBPW200H7Cz7v5GUyjz8R33VJwWh4J3rEJCeHzPggAkj4B8V1kT98fdqp3yH
9mu9LS/tEY2pl6GJe8RflwlrwT1Y/HisXZMu3ulbsb/y8no7CG3HRgyH4Nd0lzb6eeSNHrYoXq9o
AT82pQCoOs3l4XobcRL9AG9P80LGPzDdO6ThuclG+Q1bsgzMBlsEVToYyx6aAsrla5wmi6KRgk6h
OwGY91963tZcxse5Hv/n9cf/fCBGCfl6ZeDsUqC56C/gY52TvXTrUkjm7tqQR1/uHyFwAjrrwXBv
3M5zK+Ws6Z8pFms8LK0uoUHbix+znR1YNVGV2/0skmwHbx+oosuolO0/SXK8yKmHUFXptNmhfGKd
vxfEhuuW71lieU/d1S58MhNpaz1zPTbU6LhqFGJChuBE3W+//zivmELCv6fKYwpj6QIavF0+K3sg
jEMgNnM8gbB0gpDlOrA5vHdNrzH/BnQAVKWJNLaJhNEldDH7YLBNFp+vDosgxghWhUh1gieSWg+u
k/b2LdxCzg3csUOAT1VEhSxlAh83jwOhp3BuRPXEaQ6lh4PnXqHgDliKPx4wZ0Jvcz+HCbDzFyKR
YD9pQooGf2CXz//wvepSS5EPg+xjon1TNKPAhon+32/OABDnOsuyxIgbuOaS6ZOatGcuC1XCNmws
oKQmrpE9SWi72GZI4UzdZLPkVfslbOvpbpXezBDkX+S9ztn45IVHt8wuAQqerHPTXdBYpVBsbY0P
KxD14KbrNCOogxIWqkB/a7Agn8apbhK+1DK0Lnjeva5pyN+V3Ig8QfTCIzeul+EJ66vqlagyQHWs
oiARU+VurniL97WR8rd/EdJ18YhXhqhQJorfM8ONLYulM4T3Y5YW6fWh06zlanqjbfscvuZ3XXrF
U2Nxq2YkrKQY4m/5GRrEJyculrx4vntNONTiqFeDqXRd0GbG1p/oH8WZxdldXy/KkJrjGBwZp8LO
L31sbX+OStMQ4z4GiHh799jgcpsoLrIdAt2NbMRzKC9tTcOUEBj/c6KHOzFyXt0qhClcvsgFfXjg
ysOHTMUrEmdM3X2hfdoHRthQSsHKT9BQvb02d7QKVIQJ1EnRLNEYmLgnwGeIFNSuy3fZwD6ULDLm
pBPTbJk/hHOQqbS/zox9wfITayetW48loVh8xJgwxkUbueOFtxcF0ZtLXFuLf56oev43e+vlmisn
0DViZ4ldhGzAzTiY0L6UckZEuT+uJCl0C3hg7aGsWvWMBb+jnbt+8KVPsFjYe/Z1BcQ/aVz0h8j0
xIldzgzEmSNV+I5OW9L/ZrU7yx3iznEjL4+Wt7c9Zcewv/jM9Ur9WlOyidR8WZYyT/Rlk8KfRVFQ
yclNZnPP5ReRV/i17XkLhN7+9wUydQ5J3mgUqukOomQlcShTg7etr3Brp7GTUNKvpkOEEFMb/CYN
Pox9qk3sxbv1O9j5yctigm2FEUTIaybPX1oM8ixrPUvhJZgZFZ0lYhZYUiTnvpL6Hki1CnnTUMBr
gCAarfbYtbIWFkkkCYBSTvnNfHcOLfDiDqeWfQaBXEBoWS7E9Ee21YVeHUdELg/mydELzgGLJw36
hzLB3WAZCwn83LGe+agyrMlBy6a+8SNFCzTz6jd4yY1IchCXrGU4pws4c9vJ2ObkhREkcGGxm6W2
vzPFqDOAXUgElOQnsVJ2D7FwYwVmhU26YONGiaBdoJrpYN0LJ6i8+dWzby3BqPex0cM4jMR+NOOx
gqRBolwLjZpM1uDk4wiAd4Ub/N2qeDKH8dYqo1GRCDo0yniVpuUhuoTVhNFtMlwwMQwKKBRb1XId
mC4MXMfqPCydyV2WXwuK/EHVhFN+7ntSD5I85wVSjRxslV2Fk9TyvQef5k/uhqh+NzJPP/ZsS4Cs
T4IbivnwkuFXy4czI5PnWmFtsem6A5kk46JKX6Qwa5jEEBWIVPwxEe43dP8d94DxKCyl9yor+vNN
VsVZo17JWGu6Bd3oUnfCqNfKujGw3mkfPkC0m6OoI44UGbaZ9rUBz6CsfHHZNLMqxZo/MHhtmJfG
6Aro+FOK38EFL+M7G2dAmHKDpPiJsiG33vUvre01ftPDkGB/UNQIsnr8/a35INXGe+5gNmQvzwCD
HW0WdQjrPgVOG7/YuUZrmzQc5IQluGGtQ/lbmJy2e9vUdgrCkUyxs0BSILwPpgIz2Hi3+qfsc3iV
v33U7M4MNv9oB+9VE1yyJMizMQ2Yq7BZU3vRKCyGQZ6pwqUpO5XGK7aNG7+VGJLQOJ4Uk/OHP+RO
vJOyvbVosbdfmEaoDlZ/pV2/oHjkojlUO97U1t416V/l7+AR/lEgtXB05HILHZ95eEelNUU84Aq4
1Ml5swyy5i7YH+/ISkUFc5Cb5oZRH5fdIZB8FLZO7YXaP/BFcdPXNn/slL/wSTL6LWhfZSPtBIaH
nIQq0OV4K0wz+hqHs+8+Vnb+wqTy0afjLwiR5ivWakpqC9wT9SlKdLUdqZkNHzhnKN0E+azce74p
GHWYjrNwdA55V+c3Xii5Cok3Ea9Ea3UutjG3bUf3IBUsNMMRZkMmsdv3yPJsSJLEK8Sf/vj9ND+z
4XqEy+n+DL2G/1fV2t8XS5W1NEY4WAH3g1cbOgk5k+57Zvx5P+jaPUzoYtfakQG2IEfSziGSZkWc
B/W9zaAWrQ6MWjl1qKvktADXbBvMBYFMvBWBynZRZ0QhIDLfOnw2c10+lUOOagpHpY3w1BG3jDp/
L9bxzMRNAMX/Y/Z3DDH5NHpgfPgdUdICqCVVpH+dy2IRppb9i77bmnbJKUPBDCCQY50TnXZTqgjj
aKr+mBtfq+wISETqkkzxxhzdhn/g2giX1peAZXKsCudiRX9KevXhOadKDWLuhNWr/pCLMOe6ag+F
kQ0LYCK/X6000O8Qu9HWGm8fwIR6ybb6R0A277818j+w4IbYGiur2UQ9bt9419LBc9XRlGlnr12l
bHhfirUQ6IL4ebi6Z0jx7hTpN3ixKoZL+fLw/AZnhoxbJ0AOOCn1DD12XKm5vFQa6Gl745rDq8Fc
W9wRwnNwNFDma1z8ESjhvE44hJ55c4OvvlV2rYCrTt/wOIwieTusZ/Aeyz1IogeOa6dIMkjidcZx
zDq/qKGP6HoT6u4+GyTHt8JdBvk2HlJeouUJYi9Jq8d9PNNMVZzFDk/DqSd6tIzhTFj5tjEYoz7d
2GlS9MVrN948GO03RjAvjp5Yo/752cdYBI48SY81Yn2MI4vsdvnz1+w1vy4rIEGT5byRSqh0xshR
bWIVv24w41T/nfdivtp5pwemTPZcG6Yog8s3p/uEewYhFhBIL2fYjsAZf4Z48Mv3C5ugW12nvZ/i
J3ukC9H3JlABBP/imXgZarrchJF9o8Fiiam5vjeTGuiZZHlKBaCjEwckGh6T+2z4evLIHRHZIYEp
IkW9VS7uIE8uAJtdNkerdN+FASrD/PoFr/043GSLjv60N+qeQ+MLe7S778q+TDznTGgyZtrGgZ0K
h+wEyrSZnOlyQ25VbJ7DLDnKILs1VxZ+x00chBUjVm6bhldBAaEkwn60k6YIyv0Sarad0SJWmVpz
LWqcQPhXM3eyrJF5O3tl2JyASsQsND47H1T6WeTZIFLOACMwCj0RvGa0YVH831qDuKY+R1JhUT1R
BJPPmoiHe6WbC4QPP6oEaJzR8CqHh52AhBn6J0vmzu2MmpZjsJk2A9lfT35oS/IARpeRWVxl70fE
W72AWhCq3kEC2kNcxus9W3GtLhF7G+OLzVTYU0QAXfrwevaIlb5G1D+sDW3/94CGHvxrV53P220i
rTLHmhG699RN1bAuqoS6YSQBgLl1ANRXLpZ1mtpj5TIPhx4de3Q9A1FIe+R9GIjjZPmke/tVEvS2
x6mnUCf6rUHu3BHY+ZIynQUOASedweEOnWCVmyt9Cx8PLLePbN9l/UBqYNcYo1RXdAn9o0JUdOo/
z3xHiX50h2vr+BM+oeEGsMTNAxnc1ieMU1OCffKxJwbAKXhZLrcfCShCv4Lj/a79UCK4II+ItSd9
BhhxB+7wsiwPF4HNqVxKlq6YHPtOMT5jFzTSfKL6JE+yd7qg88NpMYGH1XRV1oQv0pn8WtYppLBe
Rahf4IJtMp+qGMRXP09LQi7/OOTqAUDbxMvfO41td8QM56zuhV7SfrJ+vOvOJ8CxXuASQt6lEI3i
irw4vMxz4N1AzL8aeBdEDIidtA/i9vzG+5IyGuxil9onSOFprmjcYFcWoebNBnzp00yBnke7i4Vf
iNojmsRppqTfaTi+Ns6kOILrJM1K5g4HvuZ0oJANfh1vO0NWFgcZCzTNnVb7pj5YwiTe1WMmtcH7
vn/VxRBnYrxaj/IkE0AXxPOyak4vcJF74ZnEWNQD38y/mcx9Tl9dp46qvPgoW4izIP07/ER+amvz
ziwxtYFwB/OsSSREnKFbjKVM47cemXe4NQW828R4YPRiwfOUkxBUxGCl0yTAkH+R+mWdfRhKf4AY
hvieStCLzomeGx1aVUpS+0h34HKYbRltUmK892h4j9wwim2R6BraJytJBKKvLAKc+gKdScMgB/oB
D3M5oO/P+Y+KZc16VfaAbWgB2ZzVwv552mSHo8feekA6fzwGqvBSo0psmH6apW2u4xfNRERMoXuo
vywV00gdlk4RyNW0lhwv63Kd4EPAQ8OXc5P56Q2tTy1/dJchDzrnIQ0bemulWEVI4mCw7hfAZjNi
Zoq9Ei12GDIlAz6r6ampCicv78Ef0ubcRuW0B2l7cr3Rhfk5RARHEZ2SOe68O3mUOK9r8gM+QV05
DrkdV48By/fUkx9pbVQ6DqB6iBXDG81ShORo2BzKoJP4Ez+NR3S3EzvTu8t75GX14kDmUDzLZqnx
/XdCNskKaVql4kxb2cqD1HTMeR2DA1hg33Y3Pw7wmGNluBItyJU0B6vmhhwithFJS1b1/CiuGkgB
EyVCh1jOBrkiVg8EEyTd7gK3aZk7GawaAye9qsSbFpxy1vSjC95Cz0pBjv0wi6H0DZrkQdNXdjSp
QrTJejxbfcrU9VXzSJJOSbyIkWWRaejdOnyivK0ZJqQNUxtSutcl8mQuxJ3xOfttBeJmEk1ABpsX
zqJiv7HUrRsWJdmMLZzFUup7FXwzpiWeChWZz5SntsA+f4OjcE8n+cyojl+NvVH/2YJuEPaK0Jvm
AFm+P5er/MyxBuj22xfqamZH7FlyWtSqx2VzS1nvjwmnnl7FKIxJYpMYvIj4HiGdsOf0uxUiEOjl
wirP3pe+waiBDWZ+seg36fs/ayYdR9vwwXJNiV+XM2rIpRbh6qMFK+AT2lKaAViMsh1PKjzmqzIW
bCh5z3RuZ2tRYs8R8Xz7P6bT2YKm4Xraq5S2lE7DTfAvqx/BZAg2/BHeasied4scjWFdsxrKw4g9
bzgvgg8GYkx++99Z7IOHXKUus3h43BsT0uXfmOO3MDqmo8dA4kuoi+j16ST1mx5f46LC7Rcq2rGH
JaFsFdD/amHyyeu/U1KodnCs31xwxsgj8TfXwneMYlHsYK3ZmtoUTV1Je7WFR40Lp9LfhBdf9WkF
dJe2e6TyMNsgQ6nqr9jwtxDKvEkXdrb+Crg/DlD5XLc373QIa9uDlPwWU8dyP1/Ipl9Jib+ui0em
n7rCZKkcHpvOxEzrDiX79Ie+eqCH/y3DvESkeotMBq19YQPQgbXIWkO7UfKajKYRWzpj/Dno6BEm
lyPNEQ0Hql+uKKQUJNX3HDsFKxIj+O/8f+gu+M2/rQpsWJLjs4KuZatLtRkvAi9054hG6csYU0IX
j6fh/Cx/P+NfbwzZoNhRm0pYh2zBuo69OHNBb3JZ8mAf1/4/soUQLep3FSJBC0ni1BfSWN58Hv/2
9quNW0cyLT9BLBlcXYi7CboDnw4/rNgqyULA2ViQQlWaH1GuRLSysFp7Q6wmxBsyOzT1gBEaSyEv
UR4XhsTw4/ycQC2ZlBCG7BMsrb8nBHrp37QyPQfsx7NgpFAKusXSdWKv0fhKyQ2rPCAtvzXCA00e
acZ2SdwGtrP/9b67EBUEI+F2xIeyOfkpOiv6VZU/OOPLXhXMrvat0Jq0FDIdzF1k4AQeV+DQabGk
IPSLrFTdrlWK+tu7Z8qvL187Rdd+PbRgnTX4z+RS0Z8wdLPst7VNi8AfA3wi5e3vuBNfo0i1ucKW
mehSkIaW5AF2oWAuhxt8GhvlUwamWRhGv/GfukiPI6oYFCnWZAI5eOiTzGWt0O8WWmi7kTaombPO
5qW+s3WQDSBvfWSBf7eZ+l4UcEl2dSGLWxl72hpvP35Xz9VBxHxDJBXVwmup+Zyg0kvihT8qjuDd
+NqclNNjZZq4NLsRGBGQHJW7BDcFRJDme7kI3Yfi8yEKOR/UJ+odHGydmvIiCXZcfyr7DZlhdio1
Vc3WoBz2RQ0TFfFlGD/+saw5li8BeWU28sKb9r2JwV2TXhGWML/SOix936efWjlwbyxzeYrEnHuS
1cN6qcyjo23EFVshyw+3yzqC3VWUk+5htapSNTkcTjypVNR2XMdtRtW2dPs0SzMpr79NI++oy8La
ZvO8qay+A5UDgjeQQ9UGoE15K4Idkb0YCkWUPXtZ2h3dCH3zjUd3QZXj2kvMUIZ6KlWJUfESQqgV
+uKdQvEbydnaztTxCjdJbseSyLuSXBMvpUwxZRLDmEv3APpaeMf3mbNGzzt8lYdE+jNQ6GA4JMY7
+jnqsXmCbKdKIEfT3mN3veUU7b7My1aZP7aPrRvJq1chbjaDJZybAILz2qWEeECXqqf14JXC1tV0
R/5NT4E2z6KFaL/GNfCHg7WgRR7YdfdiWgIUlVFcW0iQ0MyGJAKg+pd51gzcvsOOsTznV95aM6hc
s91GY3ZBVygjmrbIFHL7OmJ3d86NHq0bOcMU1a5mMha1C+XAQnA3AeDMiRhMYo3lcHzl/KuGgKM5
xM0/26wJGq6UHgs5WetOkKxop0jLk+isWj6lug/Uln1EX6cMem79a4jwlvpNiiGGjQKuaW4/H4dy
+Nn1rkPCqYB8MGQsSsiMLHuQls6nB5d2iiz3UTd0HvChr1OhYwZ+XozJwpUfNS5cQZKHFwkHaFNx
aIiar4JSPNWe/rpMfIDVrAz05T49hS+G3pLqumJjoboP8oXKjJn4gnOlU69MlXOz9aYOFy9Uidzr
Zao6+evgbPdbPll7LLra45riYqrGR0nPI2i9zPbmzCG5bSobRpbQteC9S+73xExA/sW1WXFbveg4
gFhZQF0ZPWW/CNQONZ8PTV0zkUBnIAuV+ct9V40QGKvBYh/yVdMF1qirGaPMxCDDBBxepCx/ceEm
/HRGKu4CXua0vcoEzaw9nAjsECo8OpeXWaeifGvGpOyL/m05vSknQHyYHbJ1v5FUTI+YunzjOYaU
p5flFItZ1Aa8+JrLZVBEVIWmmNp6PVtGrVm9xjfTQ1854odk0Y9PEtRTs6xRL1Jx7QxRZdOMJUG2
wKu3MKVa8QOivC8oOYUIQO9bBzfT17iCpmil62tcI6TlrrQIFmHwImLQPI7XVtmKkPjF1FGEDgFq
/J9Yg9MGj0HpwwRNwM4bB3+Dkg6HxsObr+lg1MVdUWruZkoVeypx/WK2eUAOvINQ9vLIR+KEEftI
7ulkH0pSwFpXsNv7IarGsxYK4MJKX6MgHCBDrjvKu0H96cyfMTy9AyjU9Q2qmTX3styuJEsyIe/c
L+FJfQDD+tovG1LhUR1jUGcJs0zvNWMvXk2Up51rnyU6hmYMn6rxSTH3vs9nRcsiqCfdX3UOVVp8
fiiCevoBDaxZ0dSVC72Ihlv6OzKcg6YTHhoiflEugtS0knC+Jaslf4Cs7/RCxLhXY2xADEd1XDmv
AYO/Xt4iG4QCTl+79z4tonsC7EB1xA157K6nma+IALyFa+c9fdboD9PyWotUSf/3DfOTsHy1TF3S
ew58z3nkQmyxugwXybnoJmguIfXe6tDe/b7g4A2KOWhhyRVgb2hsvXc3Lvv6oS9W21al/8V1CQv6
2LkTltTnlYV1iOU/fKlbxm4To58alLC59L00QpBdRr5RXrkKNI31HzY8m6o6O+WdbnIBJncqBilL
gtz/Pkmdzp4qptJpD63IyBcWcmuKuMQoqWz2M4quFTUz/IvwlzccqP2bnl6W1aL+C5osH2X7pnOX
bZDUdEBoX3dr2rfzwYQAFXshjBB9vrY0PO995IARGNGu1nR9W2YUR86Kre2iU4sn5jk2PZELOKpc
HIyLAcMeeF73uKMzdmN2cZCLmorbideyOwNShe23UaJU0CSLzrsW7xQGyoA1iGCqpjBljqU56uN4
yenex2NbU+9waKO+OJV7Xn/UeUHJ5EfYi196HcTP3oclIfI75M/HpWJlUhlBwNfQnG8bHkseuAAc
9Q87NBC54MClQb9VN6Z/gJVCTe9w+58p2q1kBk95m6ovK0XXj0ONSAbUR0meU+kqPQUTR4LBTIsL
s0F54pscK6HLFtel2UOAJLobYrXGc0Bfu73h45Q7hgxUgzi6LVLNXtqRkWojOXhHwgrLGLthlCVW
jO/LkGof5tHVNzQDb+MEOdKTxowoI+Cg3+xlAs9C28UwEyqTDx14XvpiQkp2h6YZytrt5PPK4k91
b6mEsAZX0yLx6CbrOybYLI9xY8EX2+dfEtDt0vKOq3Z3fJQluBS1UMbPJPc06iyzczwzeUXHgxBn
68GM3IFndBV/enRSzYQecHT68UTnl/fFIltNP0bGEf7RdqpQZS8PfTBs/UV2GtOv5/uZ1PQfipjg
tSBHE2rKllDPxdcS6w1D+/twYU7W3Wc56TCtZZnYK12iNd3f+V1S6Qinp2HBoUxiTbRUE/KY+FiG
Qo36w7DDrqqOvltPFp6wtbwDmdF/2ltdHaQ4Utvd0RGo8wVDhmNhxRbqioQkckkXCTRGeQU/fW/3
3xQh3FxkOKkiPM0wJ2nKBch3lm2BPufUw0jtQqpM/Kp5THnm4CyroRzyb24x7ukup47JJ+OfoBPL
rOBsWiK5O7DcZWpxO/uc2Kd1ZK4KeHPsDTslTxHhUWfaEux5T+PFKLTubvhgovXPG1I1NPnArdTc
ucVwAHUmmzRWOdBhbmxZ8JP8nqcMySVJiuj6MhMzA1GfLlms6DDat+ppAREymw2znERyQ4to021c
QDIXml67cBQDL5sFJFwrXx6NaiIvkaXq74FwgrDvGDNAQdKLBho9u33sULr5/SiuChBegC6gnfaJ
at1NcDKAnLvo/3kyycCbTrR0TzG0d1YpggsdoEceImsk7Y8NkeeMAmFxt/5z98X2oxb9Rp0GFWHM
l3+tNGCgm/Za1aSn8piMEtD7GcbXwfVZvk2q4NYnpeOQTul/FBekhDmJPG3gh952a4gIVwdxXzBd
XW8+KC9/4mjsIUQGpDJpOcRNLmEh4YTFJMAdJ1Rb6qkCB92cBNybB3oyzqARXSkHjvSA3i3GKogY
yXDfXdmVWYHOjHESksiAKKhjxxIOnwYrH+esYYhsn9ieh5CoDf7Slle+/07fiyiGnT4yFdp1jAUu
aj1iaksgCCLfXMe8O6BjxlvjMKoAuUGK6BWw8egRr1IGVP86lNivC1c7zoSvY08OOW10SBg6D/tZ
hzNB/R7yYOHFGthiXmbeO1Sbr2H/f/LsZZxEMh5kDWhaLFvKyJsuD/LMxsJU97eJqt74oRRgQOCt
E4f3mlMswcK9euGWJEJUiSYe/1ZHApu7Wni/uM2Zpw4xdsNx+NDgi25CsUgrRQSPIHTMCn0f5CBA
ykqh8jAgxa4PxxTjWbDW87dEzo3LZaBzB36b52muU0hRxA8x2Brrsz8sAilCKgKmT8vgpNUEsSSK
gTRi43ZqELZyzZMsUcRV50Z+yCgDJkBxRIV4XfCzzdYOt5y4eJlJF3lVA8qssA8MhrxSFgBnbqGD
xgwFdPf3HoxlVqK1qhVkqx3W2DF8tJCdfhhYoHcKUUYk1kmLRUBqYtov1RM39XRkfHs7v9CqyCN0
Edr5EHbX9xC+l11mfZL+HWz0d4/ig10ZltgxaPHkrrTuQF0QQcBSRrt9AHqlsXpeWLfQWEeZ9rmC
Tg/FXskzCew2YnlDmBwnsfRvdgmgR2SFs6i0n0NpFTYIu/q7m9DiMVv4kW1alQQDD/6HPWvnQ8Mw
EapL2BQamJUzF4T9bvvHWIKVSq17mT+28GiBJ6bQolfhSu5sRLU/bWjBlGKAX55L5B9FspqkOKHZ
1FbyYKjhNXqgFZYJHGSRAk8Yc64k8vug8/PRysN5nHiUFT8jo0EvBZMfOz0ipzKJ7skkxwMSZw6S
hatOKGJR5GKpxXZyOsRHtMAhiKu4rpRJPkOtmN5uxbC96X6hmqmDY24HcbvC+rkkY4XXEHn+50Un
ed/cZNxyyhu8jeQAMdl3RK+8dtDctOa9p1OZcsLv2F3YH9Jt1jiad2BHLslMxbx91hC1wZtawUgV
gQLH7PYLRP+llY+7+J1YiC1G7z4xXCM5PcVjDMLkSyB1hRQ+NGj2vbQdYpYwDSfIprbXbpMWKzsW
0smS7TsjGeNp1sg7EoMR5/GwOKig+eWTJDNR4pPDuQiTKjq7x8I9uie7PGLnfJCzwsczHGzKNDh3
1zlJ9vUHkhOug9P3jP4PrwTKk2ax/AnkDB+PrtwLagub3hQFF/lPNqRJyYgksVMTQb+Q1f4s+cqa
PV8eSOC7E4EsNm7kT3milT4WAU6bs8Qj4h4DS7u0k8Fxoa8M9hd3ipqCEBaZXbyCfx1Rd+zpn4u1
Q1Xq1fCOFhYHxHKppnafpqo+bxxaWIkI24RXCq+9Zn5XbukMsgaUgMi5A+mLh+GrlMGlyJe5QqZT
HVJF4fJwqN4dtuiY7DSPL2MFudw3xg3qMtFMQoZsdLALnsWWcaz1kSUBFLsWqA90yKf7wPpgm3js
TFMkQXbAckebNBqkVZOWzTMl0aVGExL4kadodQuEJEUv3izQFTc/QhrUBbl7+WEpIn7ZyNZ90PKg
lovBZNI+qxZl3VikEdRdIC9JUguGhUEl2+O267eIhCqeiYhSLsalEgq+hp2aajERsJqwWYeyK0Gr
SEay7oVJXA6B+VpF6xiZjYoVxWN5C8dUCVk4hFpwRY7GhvISdm8SQWcZm7d6wyXAWHhVXmiMWaqD
aTEXj36dFPVKFBYzVehKezROtdKQReXYBcCi/MshR2bpZTf8/XAWwUd9E1XbStIhsk9W3OCVjZFa
+BXZ5yG7moAC8PO0vPpOD8P++JCR1ydIDlF0C4v2fhXciRkt97GdwHNxtMyzqEALEnicifTjrUo/
U79t9dcQ/w+ChiDO0LO4fr86vDoV5YDASHkorF6yrtrawZv/TtNdNtbDc+tOMeCQb54Z1ByeSeRh
JPOSjS7Ki0Wjq9YHiCSjFFmgUgOGlLYc1nXaOO6KzceLwM0KmGb/wOvETZq2+g6EKT2mWVSoZvgc
VoYpvVws2eP8wRIqapDI/eEaQomIiPjBemjmwJ/seA+R0D3JTNmY8i//31iageEfaiUQ39S2e7bn
XynmgomS3YIgoYFDpGpstH2oC4MCv0ezDP1/3JfGjC3I7PzHFGh/wq09Dn2347gEjSuBwavykPL1
UzA68hFFl3AdS1+kinc75UBFOj4E3l3faz8E/yIkQHcavgGhInPv0Iv1gkLdsHIYfK+J8cnGzcKi
qWcvnvVmGSTheOK7qPs4b2z4LwbKa0bMfjsH7uF5v+y91B3j+BfMbTj5EOo7WUBb2dwxPpgmcr3L
DxcJZqr6N4D5Ihm4Unt/8igwIv8vkLIcY0SEXLwdshjISZeGnlnNrxMJV2+qp1TFDevpFAOVM0kz
z3cHnf5JMquzbKVgRwz2gtKz7SPLyA0fV+tOtCc+LOuLQlK+2ovNBCFICnZaI/62/NBlKfo2Hnz2
sIt5F6lWz/BvWMLOmOrrQBQto2u11B8AY5NSEjs3TzcczZtXobUgM4Ph3AFxjKss+KQdXPox0MU4
kdMvYLj2eVJdDyQizMSy1aaSOOaK5pZLFIy39SFhOGnec+IXltXSn1mFyZIiwNa0kH/yxLO7MIW3
AjuqBcVOvQAklV01MwPjRhwJvqiGEh8414Pf2ygSbeAkrHn+owXBt0FaNrTxi7Sy4O+CTSH1BREk
t8fRXqSnid03Mwf8qUli0eDDiGmVj3/aRJJ+C2hpka4CJ1pzokncK6NguG6R5bR88KG6fmudgBRA
OIFoecvRIWHLTwQHZuXbZnItUkmB2UVmML9ie80V04YPEe5IYlrmDkonJdk5pjttP6+1KUW/milk
MSExUq0Z2pu2MeNmF/qzzrpfcb/I5rZCMh3U6x4hJVZgw2Y2hL/CHEWIAjq3Vo9pwSj4cHQGfsNn
q9yDUwiggUfIeqgnec9u22UPe4MkLSJV+Kk2elIPjxMoQOxZ0nkp1A38uTIHA5LQc8OIOD1tNFiL
cwGU3uNw5cxuNxIYdMXzwypUbCYaQ2LLORj17c4Tz/YL3pm/tpEuphCIsqK7//Z1I33k3MRxUKYV
lmLIGKaf7WKsv1YM9hLuJku/uJ7iDsHos23REJ00XWiEfTa8LnJJVNT8ILQ0gXUTdjTmHunFvSAI
e1q6mTEn1FWAHfwG2Ut18HQ+Asa+F5SDZA/P7T32FjYQ75mZ4CXwQCYJZymidOCRFjJET20+xdhG
FGHJJe9kvElip+6G0IpGl3Njj+ol0y6Hj/vM5j5RCLMS8Eyi3GouzftdA60Vfk7ty2Yulr4dBMiF
iigXT3lxAjRaJ98tSUG7ILYju98iLXGL2oUp3cOsS4bTbwEk17pvdRpqoBMKWatOD82xXp+B5yE8
y/ngt204fMOvyFzDqCpeEZufKR0BvlG7pI+ggXJvF2N+qazSwvrnYatZLOtlQAxUrSxSaHx0LMdh
CI34cBGYIAu1rmGGnIJDNzrs1SQkGdtaBr55eP4OZC7ke0uLAmUd4ts4EC1br4xFBOxhW8UIl17m
14rJMBvPlwe9HysiXc0tKHI+1j+I2eiZdHKkBKEAo9umoNmGznJH+WaRP70LKZaxzZvfiJAkRjDR
SoFQG8/G5WD2r3XJ2aAwNdhkLprR1XLzGyDnemtYvk0r9y6F/uHgTdgYg1MS5uBbvvLPeRWGYNOg
AhurmaQI7iZ2nxtf5pf3J1JA0xFpeg7HAEdW2wPvozjq0wsqhIzqxZPwvpRyd9DzPm7zo2/KW5hH
y0wBSNy7W0ClX0/ekDbvQBOZXASFHe00bZyevcjE/RXuMajyJS2psChJTVWnbsKhs7ihnLu8k5cP
7STe8eq0IvfyXEzcQIdggT3rq3MIQVrjTUAsylBHBFud22tHD5i1do/btetbGCuBLxYieNh7ccrq
fdZj/NdJ90eekbROFf4Ai0p5u8grE5hApy6/F4Vr02Y81Hife9lmGEniST1GNstKFdJrhYCLyY/O
yWnxZlEjQrV/8txghKSzQ8PV/sdb8YzhmQbUiz4Nx+d7yXADOn5XH4j9+HLq+qS69QMjCIboR13e
GCklafgHmW9ISOTT3vVmWtJDPAZD+4nACvlKlo28V6wwMuM77iPqMrOkV3HzKD9n+2a4iLTOMu5E
VDWnQd7o0g22bVK/TtYVYrKqorUHI1LQAWOn5jNhIDWdiPPpomPWqu/tGQsmyXJj2Q7CgFSQFfQu
Sj+idb++uszSoZrqhDvPgxP//rcGb187XcecS/s1vGxU3CfozVVVdJ18M9JssIjoXLuLrrKpcPgb
/cU5Pj026oHeujfHjKzqqNfW/7si6jVfkVNi7lCCY20lf2qYQ5S4+LxcYDDJbqWcSqyfDeM5hTDH
g9FuH5tkdVzU3Bc669pDc2Y6MIcm8V2KseulBN18Z8ZsO4PT/HjtQoVnaz+vCwNMZZQS/LjmRfoZ
oG7liu0+swnapU/bt2YqeqGXTwOC+kLN5PaCqKsAEDWr80ygZP4ESCO7uXp0MF55oAUn3TSA/ube
EBQkXllhBYdn2VkUyujtBJTMRMjwyn35c6UNMt1EtRlkcCKZ6r8kfKrB5eaRRA8JHoaZyMMWPS4b
0iKCWSmrhNdJyx2ElJWXtZnc548k1MUunhS28kRvbFdqVMhmxGbK4kLAO1RvLd49ho7qZcIODqPx
74G6RLtr1FwiVINySKOOYeoxIph03BDj/r8sTXnJm/yPbeG8RD+8V5uv53MkfZNiMh3txN+va0zs
lzczODfzEEkUTej4Uh5FA8c6aQ23/h5P78NGcKz7itmGxVfEm7txYVuO6pMW44Pvx6ObXdzwhnaG
V8NlJV20340DR3PM515hQx/+UWG2mqPIWCkNAeC0Asr9kIfuN6IRvcZ/RisIDBQCBsFsnKbE2puj
a5EtXOf22ANWk0Svm4e3tFR5hBtjKSkSMjmTSnancODaerF2Mjg5VlgJILjKPLUjvVqKHtGxqClM
z/aIrMhmuepUUquzRbeZlKvHh6AzMVmBl/u21rszr5+j8aDToGbB69G285xpb4hq5i14TuEcR4Ri
EDsODfqAPP8ExQdsmX9E0MxsJ8WZ7uHI1gvpmvWrQGPY6twNlhGhzD8LLU5eIDM2SDc17Hcv85OX
twpZq7tXcrZsW57MgPlRknCGKiM1INsXYSpIiEznSyKV3ugajuGil0MkL0NLST/Z7xhL4k+boO0i
RIoM0CvGh+VvMgSz9LD3pROC1GdQo/FHBQ+uJQnxLb+cZbp0BJ9mz0DTxeAf1UnWso/Dlt/Qx15C
3Q0YnkR/grPcUNMQ/JwUcf8VSwQKiphCAwIYwmTX94FAYjrkggms7ZQnJYlgpZ7hYrvUzqehu1pG
9ZsQhbqNY8Lsw2pdC2Bbfm64T6w+XmpQu8k1PeJP9llUMz8cQSZR/Dc/nbqpX7He
`pragma protect end_protected
