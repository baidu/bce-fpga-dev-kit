   // AXI Master AW channel
   output [ADDR_WIDTH-1:0]  M_AXI_araddr,
   output [1:0]             M_AXI_arburst,
   output [3:0]             M_AXI_arcache,
   output [ID_WIDTH-1:0]    M_AXI_arid,
   output [7:0]             M_AXI_arlen,
   output                   M_AXI_arlock,
   output [2:0]             M_AXI_arprot,
   output [3:0]             M_AXI_arqos,
   output [3:0]             M_AXI_arregion,
   input                    M_AXI_arready,
   output [2:0]             M_AXI_arsize,
   output                   M_AXI_arvalid,
   // AXI Master AR channel
   output [ADDR_WIDTH-1:0]  M_AXI_awaddr,
   output [1:0]             M_AXI_awburst,
   output [3:0]             M_AXI_awcache,
   output [ID_WIDTH-1:0]    M_AXI_awid,
   output [7:0]             M_AXI_awlen,
   output                   M_AXI_awlock,
   output [2:0]             M_AXI_awprot,
   output [3:0]             M_AXI_awqos,
   output [3:0]             M_AXI_awregion,
   input                    M_AXI_awready,
   output [2:0]             M_AXI_awsize,
   output                   M_AXI_awvalid,
   // AXI Master B channel
   input  [ID_WIDTH-1:0]    M_AXI_bid,
   output                   M_AXI_bready,
   input  [1:0]             M_AXI_bresp,
   input                    M_AXI_bvalid,
   // AXI Master R channel
   input  [DATA_WIDTH-1:0]  M_AXI_rdata,
   input  [ID_WIDTH-1:0]    M_AXI_rid,
   input                    M_AXI_rlast,
   output                   M_AXI_rready,
   input  [1:0]             M_AXI_rresp,
   input                    M_AXI_rvalid,
   // AXI Master W channel
   output [DATA_WIDTH-1:0]  M_AXI_wdata,
   output                   M_AXI_wlast,
   input                    M_AXI_wready,
   output [MASK_WIDTH-1:0]  M_AXI_wstrb,
   output                   M_AXI_wvalid,
