`define USE_NO_DDR 1
