`define APP_DDR 1
