   `ifdef USE_DDR4_C0
   output[30:0]    C0_DDR4_M_AXI_araddr,
   output[1:0]     C0_DDR4_M_AXI_arburst,
   output[3:0]     C0_DDR4_M_AXI_arcache,
   output[0:0]     C0_DDR4_M_AXI_arid,
   output[7:0]     C0_DDR4_M_AXI_arlen,
   output[0:0]     C0_DDR4_M_AXI_arlock,
   output[2:0]     C0_DDR4_M_AXI_arprot,
   output[3:0]     C0_DDR4_M_AXI_arqos,
   output[3:0]     C0_DDR4_M_AXI_arregion,
   input           C0_DDR4_M_AXI_arready,
   output[2:0]     C0_DDR4_M_AXI_arsize,
   output          C0_DDR4_M_AXI_arvalid,
   output[30:0]    C0_DDR4_M_AXI_awaddr,
   output[1:0]     C0_DDR4_M_AXI_awburst,
   output[3:0]     C0_DDR4_M_AXI_awcache,
   output[0:0]     C0_DDR4_M_AXI_awid,
   output[7:0]     C0_DDR4_M_AXI_awlen,
   output[0:0]     C0_DDR4_M_AXI_awlock,
   output[2:0]     C0_DDR4_M_AXI_awprot,
   output[3:0]     C0_DDR4_M_AXI_awqos,
   output[3:0]     C0_DDR4_M_AXI_awregion,
   input           C0_DDR4_M_AXI_awready,
   output[2:0]     C0_DDR4_M_AXI_awsize,
   output          C0_DDR4_M_AXI_awvalid,
   input  [0:0]    C0_DDR4_M_AXI_bid,
   output          C0_DDR4_M_AXI_bready,
   input  [1:0]    C0_DDR4_M_AXI_bresp,
   input           C0_DDR4_M_AXI_bvalid,
   input  [511:0]  C0_DDR4_M_AXI_rdata,
   input  [0:0]    C0_DDR4_M_AXI_rid,
   input           C0_DDR4_M_AXI_rlast,
   output          C0_DDR4_M_AXI_rready,
   input  [1:0]    C0_DDR4_M_AXI_rresp,
   input           C0_DDR4_M_AXI_rvalid,
   output[511:0]   C0_DDR4_M_AXI_wdata,
   output          C0_DDR4_M_AXI_wlast,
   input           C0_DDR4_M_AXI_wready,
   output[63:0]    C0_DDR4_M_AXI_wstrb,
   output          C0_DDR4_M_AXI_wvalid,

   input           c0_ddr4_ui_clk,
   input           c0_ddr4_ui_clk_sync_rst,
   input           c0_init_calib_complete,
   input           c0_ddr4_interrupt,
   `endif

   `ifdef USE_DDR4_C1
   output[30:0]    C1_DDR4_M_AXI_araddr,
   output[1:0]     C1_DDR4_M_AXI_arburst,
   output[3:0]     C1_DDR4_M_AXI_arcache,
   output[0:0]     C1_DDR4_M_AXI_arid,
   output[7:0]     C1_DDR4_M_AXI_arlen,
   output[0:0]     C1_DDR4_M_AXI_arlock,
   output[2:0]     C1_DDR4_M_AXI_arprot,
   output[3:0]     C1_DDR4_M_AXI_arqos,
   output[3:0]     C1_DDR4_M_AXI_arregion,
   input           C1_DDR4_M_AXI_arready,
   output[2:0]     C1_DDR4_M_AXI_arsize,
   output          C1_DDR4_M_AXI_arvalid,
   output[30:0]    C1_DDR4_M_AXI_awaddr,
   output[1:0]     C1_DDR4_M_AXI_awburst,
   output[3:0]     C1_DDR4_M_AXI_awcache,
   output[0:0]     C1_DDR4_M_AXI_awid,
   output[7:0]     C1_DDR4_M_AXI_awlen,
   output[0:0]     C1_DDR4_M_AXI_awlock,
   output[2:0]     C1_DDR4_M_AXI_awprot,
   output[3:0]     C1_DDR4_M_AXI_awqos,
   output[3:0]     C1_DDR4_M_AXI_awregion,
   input           C1_DDR4_M_AXI_awready,
   output[2:0]     C1_DDR4_M_AXI_awsize,
   output          C1_DDR4_M_AXI_awvalid,
   input  [0:0]    C1_DDR4_M_AXI_bid,
   output          C1_DDR4_M_AXI_bready,
   input  [1:0]    C1_DDR4_M_AXI_bresp,
   input           C1_DDR4_M_AXI_bvalid,
   input  [511:0]  C1_DDR4_M_AXI_rdata,
   input  [0:0]    C1_DDR4_M_AXI_rid,
   input           C1_DDR4_M_AXI_rlast,
   output          C1_DDR4_M_AXI_rready,
   input  [1:0]    C1_DDR4_M_AXI_rresp,
   input           C1_DDR4_M_AXI_rvalid,
   output[511:0]   C1_DDR4_M_AXI_wdata,
   output          C1_DDR4_M_AXI_wlast,
   input           C1_DDR4_M_AXI_wready,
   output[63:0]    C1_DDR4_M_AXI_wstrb,
   output          C1_DDR4_M_AXI_wvalid,

   input           c1_ddr4_ui_clk,
   input           c1_ddr4_ui_clk_sync_rst,
   input           c1_init_calib_complete,
   input           c1_ddr4_interrupt,
   `endif

   `ifdef USE_DDR4_C2
   output[30:0]    C2_DDR4_M_AXI_araddr,
   output[1:0]     C2_DDR4_M_AXI_arburst,
   output[3:0]     C2_DDR4_M_AXI_arcache,
   output[0:0]     C2_DDR4_M_AXI_arid,
   output[7:0]     C2_DDR4_M_AXI_arlen,
   output[0:0]     C2_DDR4_M_AXI_arlock,
   output[2:0]     C2_DDR4_M_AXI_arprot,
   output[3:0]     C2_DDR4_M_AXI_arqos,
   output[3:0]     C2_DDR4_M_AXI_arregion,
   input           C2_DDR4_M_AXI_arready,
   output[2:0]     C2_DDR4_M_AXI_arsize,
   output          C2_DDR4_M_AXI_arvalid,
   output[30:0]    C2_DDR4_M_AXI_awaddr,
   output[1:0]     C2_DDR4_M_AXI_awburst,
   output[3:0]     C2_DDR4_M_AXI_awcache,
   output[0:0]     C2_DDR4_M_AXI_awid,
   output[7:0]     C2_DDR4_M_AXI_awlen,
   output[0:0]     C2_DDR4_M_AXI_awlock,
   output[2:0]     C2_DDR4_M_AXI_awprot,
   output[3:0]     C2_DDR4_M_AXI_awqos,
   output[3:0]     C2_DDR4_M_AXI_awregion,
   input           C2_DDR4_M_AXI_awready,
   output[2:0]     C2_DDR4_M_AXI_awsize,
   output          C2_DDR4_M_AXI_awvalid,
   input  [0:0]    C2_DDR4_M_AXI_bid,
   output          C2_DDR4_M_AXI_bready,
   input  [1:0]    C2_DDR4_M_AXI_bresp,
   input           C2_DDR4_M_AXI_bvalid,
   input  [511:0]  C2_DDR4_M_AXI_rdata,
   input  [0:0]    C2_DDR4_M_AXI_rid,
   input           C2_DDR4_M_AXI_rlast,
   output          C2_DDR4_M_AXI_rready,
   input  [1:0]    C2_DDR4_M_AXI_rresp,
   input           C2_DDR4_M_AXI_rvalid,
   output[511:0]   C2_DDR4_M_AXI_wdata,
   output          C2_DDR4_M_AXI_wlast,
   input           C2_DDR4_M_AXI_wready,
   output[63:0]    C2_DDR4_M_AXI_wstrb,
   output          C2_DDR4_M_AXI_wvalid,

   input           c2_ddr4_ui_clk,
   input           c2_ddr4_ui_clk_sync_rst,
   input           c2_init_calib_complete,
   input           c2_ddr4_interrupt,
   `endif

   `ifdef USE_DDR4_C3
   output[30:0]    C3_DDR4_M_AXI_araddr,
   output[1:0]     C3_DDR4_M_AXI_arburst,
   output[3:0]     C3_DDR4_M_AXI_arcache,
   output[0:0]     C3_DDR4_M_AXI_arid,
   output[7:0]     C3_DDR4_M_AXI_arlen,
   output[0:0]     C3_DDR4_M_AXI_arlock,
   output[2:0]     C3_DDR4_M_AXI_arprot,
   output[3:0]     C3_DDR4_M_AXI_arqos,
   output[3:0]     C3_DDR4_M_AXI_arregion,
   input           C3_DDR4_M_AXI_arready,
   output[2:0]     C3_DDR4_M_AXI_arsize,
   output          C3_DDR4_M_AXI_arvalid,
   output[30:0]    C3_DDR4_M_AXI_awaddr,
   output[1:0]     C3_DDR4_M_AXI_awburst,
   output[3:0]     C3_DDR4_M_AXI_awcache,
   output[0:0]     C3_DDR4_M_AXI_awid,
   output[7:0]     C3_DDR4_M_AXI_awlen,
   output[0:0]     C3_DDR4_M_AXI_awlock,
   output[2:0]     C3_DDR4_M_AXI_awprot,
   output[3:0]     C3_DDR4_M_AXI_awqos,
   output[3:0]     C3_DDR4_M_AXI_awregion,
   input           C3_DDR4_M_AXI_awready,
   output[2:0]     C3_DDR4_M_AXI_awsize,
   output          C3_DDR4_M_AXI_awvalid,
   input  [0:0]    C3_DDR4_M_AXI_bid,
   output          C3_DDR4_M_AXI_bready,
   input  [1:0]    C3_DDR4_M_AXI_bresp,
   input           C3_DDR4_M_AXI_bvalid,
   input  [511:0]  C3_DDR4_M_AXI_rdata,
   input  [0:0]    C3_DDR4_M_AXI_rid,
   input           C3_DDR4_M_AXI_rlast,
   output          C3_DDR4_M_AXI_rready,
   input  [1:0]    C3_DDR4_M_AXI_rresp,
   input           C3_DDR4_M_AXI_rvalid,
   output[511:0]   C3_DDR4_M_AXI_wdata,
   output          C3_DDR4_M_AXI_wlast,
   input           C3_DDR4_M_AXI_wready,
   output[63:0]    C3_DDR4_M_AXI_wstrb,
   output          C3_DDR4_M_AXI_wvalid,

   input           c3_ddr4_ui_clk,
   input           c3_ddr4_ui_clk_sync_rst,
   input           c3_init_calib_complete,
   input           c3_ddr4_interrupt,
   `endif
