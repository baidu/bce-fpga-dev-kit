`define USE_DDR 1
`define USE_DDR4_C0 1
`define USE_DDR4_C1 1
`define USE_DDR4_C2 1
`define USE_DDR4_C3 1
`define RP_AXI_MASTER 1
`define AXI_DDR 1
