   `ifdef USE_DDR4_C0
   input           c0_ddr4_app_correct_en_i,
   output [51:0]   c0_ddr4_ecc_err_addr,
   output [7:0]    c0_ddr4_ecc_single,
   output [7:0]    c0_ddr4_ecc_multiple,

   input  [27:0]   c0_ddr4_app_addr,
   input  [2:0]    c0_ddr4_app_cmd,
   input           c0_ddr4_app_en,
   input           c0_ddr4_app_hi_pri,
   input  [511:0]  c0_ddr4_app_wdf_data,
   input           c0_ddr4_app_wdf_end,
   input  [63:0]   c0_ddr4_app_wdf_mask,
   input           c0_ddr4_app_wdf_wren,
   output [511:0]  c0_ddr4_app_rd_data,
   output          c0_ddr4_app_rd_data_end,
   output          c0_ddr4_app_rd_data_valid,
   output          c0_ddr4_app_rdy,
   output          c0_ddr4_app_wdf_rdy,
   output          c0_dbg_clk,
   output [511:0]  c0_dbg_bus,
   output          c0_ddr4_ui_clk,
   output          c0_ddr4_ui_clk_sync_rst,
   output          c0_init_calib_complete,
   `endif

   `ifdef USE_DDR4_C1
   input           c1_ddr4_app_correct_en_i,
   output [51:0]   c1_ddr4_ecc_err_addr,
   output [7:0]    c1_ddr4_ecc_single,
   output [7:0]    c1_ddr4_ecc_multiple,

   input  [27:0]   c1_ddr4_app_addr,
   input  [2:0]    c1_ddr4_app_cmd,
   input           c1_ddr4_app_en,
   input           c1_ddr4_app_hi_pri,
   input  [511:0]  c1_ddr4_app_wdf_data,
   input           c1_ddr4_app_wdf_end,
   input  [63:0]   c1_ddr4_app_wdf_mask,
   input           c1_ddr4_app_wdf_wren,
   output [511:0]  c1_ddr4_app_rd_data,
   output          c1_ddr4_app_rd_data_end,
   output          c1_ddr4_app_rd_data_valid,
   output          c1_ddr4_app_rdy,
   output          c1_ddr4_app_wdf_rdy,
   output          c1_dbg_clk,
   output [511:0]  c1_dbg_bus,
   output          c1_ddr4_ui_clk,
   output          c1_ddr4_ui_clk_sync_rst,
   output          c1_init_calib_complete,
   `endif

   `ifdef USE_DDR4_C2
   input           c2_ddr4_app_correct_en_i,
   output [51:0]   c2_ddr4_ecc_err_addr,
   output [7:0]    c2_ddr4_ecc_single,
   output [7:0]    c2_ddr4_ecc_multiple,

   input  [27:0]   c2_ddr4_app_addr,
   input  [2:0]    c2_ddr4_app_cmd,
   input           c2_ddr4_app_en,
   input           c2_ddr4_app_hi_pri,
   input  [511:0]  c2_ddr4_app_wdf_data,
   input           c2_ddr4_app_wdf_end,
   input  [63:0]   c2_ddr4_app_wdf_mask,
   input           c2_ddr4_app_wdf_wren,
   output [511:0]  c2_ddr4_app_rd_data,
   output          c2_ddr4_app_rd_data_end,
   output          c2_ddr4_app_rd_data_valid,
   output          c2_ddr4_app_rdy,
   output          c2_ddr4_app_wdf_rdy,
   output          c2_dbg_clk,
   output [511:0]  c2_dbg_bus,
   output          c2_ddr4_ui_clk,
   output          c2_ddr4_ui_clk_sync_rst,
   output          c2_init_calib_complete,
   `endif

   `ifdef USE_DDR4_C3
   input           c3_ddr4_app_correct_en_i,
   output [51:0]   c3_ddr4_ecc_err_addr,
   output [7:0]    c3_ddr4_ecc_single,
   output [7:0]    c3_ddr4_ecc_multiple,

   input  [27:0]   c3_ddr4_app_addr,
   input  [2:0]    c3_ddr4_app_cmd,
   input           c3_ddr4_app_en,
   input           c3_ddr4_app_hi_pri,
   input  [511:0]  c3_ddr4_app_wdf_data,
   input           c3_ddr4_app_wdf_end,
   input  [63:0]   c3_ddr4_app_wdf_mask,
   input           c3_ddr4_app_wdf_wren,
   output [511:0]  c3_ddr4_app_rd_data,
   output          c3_ddr4_app_rd_data_end,
   output          c3_ddr4_app_rd_data_valid,
   output          c3_ddr4_app_rdy,
   output          c3_ddr4_app_wdf_rdy,
   output          c3_dbg_clk,
   output [511:0]  c3_dbg_bus,
   output          c3_ddr4_ui_clk,
   output          c3_ddr4_ui_clk_sync_rst,
   output          c3_init_calib_complete,
   `endif
