   `ifdef USE_DDR4_C0
   output          c0_ddr4_app_correct_en_i,
   input  [51:0]   c0_ddr4_ecc_err_addr,
   input  [7:0]    c0_ddr4_ecc_single,
   input  [7:0]    c0_ddr4_ecc_multiple,

   output [27:0]   c0_ddr4_app_addr,
   output [2:0]    c0_ddr4_app_cmd,
   output          c0_ddr4_app_en,
   output          c0_ddr4_app_hi_pri,
   output [511:0]  c0_ddr4_app_wdf_data,
   output          c0_ddr4_app_wdf_end,
   output [63:0]   c0_ddr4_app_wdf_mask,
   output          c0_ddr4_app_wdf_wren,
   input  [511:0]  c0_ddr4_app_rd_data,
   input           c0_ddr4_app_rd_data_end,
   input           c0_ddr4_app_rd_data_valid,
   input           c0_ddr4_app_rdy,
   input           c0_ddr4_app_wdf_rdy,
   input           c0_dbg_clk,
   input  [511:0]  c0_dbg_bus,
   input           c0_ddr4_ui_clk,
   input           c0_ddr4_ui_clk_sync_rst,
   input           c0_init_calib_complete,
   `endif

   `ifdef USE_DDR4_C1
   output          c1_ddr4_app_correct_en_i,
   input  [51:0]   c1_ddr4_ecc_err_addr,
   input  [7:0]    c1_ddr4_ecc_single,
   input  [7:0]    c1_ddr4_ecc_multiple,

   output [27:0]   c1_ddr4_app_addr,
   output [2:0]    c1_ddr4_app_cmd,
   output          c1_ddr4_app_en,
   output          c1_ddr4_app_hi_pri,
   output [511:0]  c1_ddr4_app_wdf_data,
   output          c1_ddr4_app_wdf_end,
   output [63:0]   c1_ddr4_app_wdf_mask,
   output          c1_ddr4_app_wdf_wren,
   input  [511:0]  c1_ddr4_app_rd_data,
   input           c1_ddr4_app_rd_data_end,
   input           c1_ddr4_app_rd_data_valid,
   input           c1_ddr4_app_rdy,
   input           c1_ddr4_app_wdf_rdy,
   input           c1_dbg_clk,
   input  [511:0]  c1_dbg_bus,
   input           c1_ddr4_ui_clk,
   input           c1_ddr4_ui_clk_sync_rst,
   input           c1_init_calib_complete,
   `endif

   `ifdef USE_DDR4_C2
   output          c2_ddr4_app_correct_en_i,
   input  [51:0]   c2_ddr4_ecc_err_addr,
   input  [7:0]    c2_ddr4_ecc_single,
   input  [7:0]    c2_ddr4_ecc_multiple,

   output [27:0]   c2_ddr4_app_addr,
   output [2:0]    c2_ddr4_app_cmd,
   output          c2_ddr4_app_en,
   output          c2_ddr4_app_hi_pri,
   output [511:0]  c2_ddr4_app_wdf_data,
   output          c2_ddr4_app_wdf_end,
   output [63:0]   c2_ddr4_app_wdf_mask,
   output          c2_ddr4_app_wdf_wren,
   input  [511:0]  c2_ddr4_app_rd_data,
   input           c2_ddr4_app_rd_data_end,
   input           c2_ddr4_app_rd_data_valid,
   input           c2_ddr4_app_rdy,
   input           c2_ddr4_app_wdf_rdy,
   input           c2_dbg_clk,
   input  [511:0]  c2_dbg_bus,
   input           c2_ddr4_ui_clk,
   input           c2_ddr4_ui_clk_sync_rst,
   input           c2_init_calib_complete,
   `endif

   `ifdef USE_DDR4_C3
   output          c3_ddr4_app_correct_en_i,
   input  [51:0]   c3_ddr4_ecc_err_addr,
   input  [7:0]    c3_ddr4_ecc_single,
   input  [7:0]    c3_ddr4_ecc_multiple,

   output [27:0]   c3_ddr4_app_addr,
   output [2:0]    c3_ddr4_app_cmd,
   output          c3_ddr4_app_en,
   output          c3_ddr4_app_hi_pri,
   output [511:0]  c3_ddr4_app_wdf_data,
   output          c3_ddr4_app_wdf_end,
   output [63:0]   c3_ddr4_app_wdf_mask,
   output          c3_ddr4_app_wdf_wren,
   input  [511:0]  c3_ddr4_app_rd_data,
   input           c3_ddr4_app_rd_data_end,
   input           c3_ddr4_app_rd_data_valid,
   input           c3_ddr4_app_rdy,
   input           c3_ddr4_app_wdf_rdy,
   input           c3_dbg_clk,
   input  [511:0]  c3_dbg_bus,
   input           c3_ddr4_ui_clk,
   input           c3_ddr4_ui_clk_sync_rst,
   input           c3_init_calib_complete,
   `endif
