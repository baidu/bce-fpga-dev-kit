   `ifdef USE_DDR4_C0
   output         C0_DDR4_act_n,
   output [16:0]  C0_DDR4_adr,
   output [1:0]   C0_DDR4_ba,
   output [0:0]   C0_DDR4_bg,
   output [0:0]   C0_DDR4_ck_c,
   output [0:0]   C0_DDR4_cke,
   output [0:0]   C0_DDR4_cs_n,
   inout [8:0]    C0_DDR4_dm_n,
   inout [71:0]   C0_DDR4_dq,
   inout [8:0]    C0_DDR4_dqs_c,
   output [0:0]   C0_DDR4_odt,
   output         C0_DDR4_reset_n,
   input          C0_SYS_CLK_clk_n,
   input          C0_SYS_CLK_clk_p,
   output [0:0]   C0_DDR4_ck_t,
   inout [8:0]    C0_DDR4_dqs_t,
   `endif

   `ifdef USE_DDR4_C1
   output         C1_DDR4_act_n,
   output [16:0]  C1_DDR4_adr,
   output [1:0]   C1_DDR4_ba,
   output [0:0]   C1_DDR4_bg,
   output [0:0]   C1_DDR4_ck_c,
   output [0:0]   C1_DDR4_cke,
   output [0:0]   C1_DDR4_cs_n,
   inout [8:0]    C1_DDR4_dm_n,
   inout [71:0]   C1_DDR4_dq,
   inout [8:0]    C1_DDR4_dqs_c,
   output [0:0]   C1_DDR4_odt,
   output         C1_DDR4_reset_n,
   input          C1_SYS_CLK_clk_n,
   input          C1_SYS_CLK_clk_p,
   output [0:0]   C1_DDR4_ck_t,
   inout [8:0]    C1_DDR4_dqs_t,
   `endif

   `ifdef USE_DDR4_C2
   output         C2_DDR4_act_n,
   output [16:0]  C2_DDR4_adr,
   output [1:0]   C2_DDR4_ba,
   output [0:0]   C2_DDR4_bg,
   output [0:0]   C2_DDR4_ck_c,
   output [0:0]   C2_DDR4_cke,
   output [0:0]   C2_DDR4_cs_n,
   inout [8:0]    C2_DDR4_dm_n,
   inout [71:0]   C2_DDR4_dq,
   inout [8:0]    C2_DDR4_dqs_c,
   output [0:0]   C2_DDR4_odt,
   output         C2_DDR4_reset_n,
   input          C2_SYS_CLK_clk_n,
   input          C2_SYS_CLK_clk_p,
   output [0:0]   C2_DDR4_ck_t,
   inout [8:0]    C2_DDR4_dqs_t,
   `endif

   `ifdef USE_DDR4_C3
   output         C3_DDR4_act_n,
   output [16:0]  C3_DDR4_adr,
   output [1:0]   C3_DDR4_ba,
   output [0:0]   C3_DDR4_bg,
   output [0:0]   C3_DDR4_ck_c,
   output [0:0]   C3_DDR4_cke,
   output [0:0]   C3_DDR4_cs_n,
   inout [8:0]    C3_DDR4_dm_n,
   inout [71:0]   C3_DDR4_dq,
   inout [8:0]    C3_DDR4_dqs_c,
   output [0:0]   C3_DDR4_odt,
   output         C3_DDR4_reset_n,
   input          C3_SYS_CLK_clk_n,
   input          C3_SYS_CLK_clk_p,
   output [0:0]   C3_DDR4_ck_t,
   inout [8:0]    C3_DDR4_dqs_t,
   `endif
