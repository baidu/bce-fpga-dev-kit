`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
U5Gk7fay92T1+/rPL9dkXOzFS9mYB1gmErtGq1hGh2NDOhMhsap7zWTE1xOE2L7oOnHip7QnOqgm
f9QlT0eOSg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nDm6XgdMQfJdJ/uDSKHMaWqz/MQCgtZ2iNjW8+CwJ/U9MGWdsBRx3ijlNS1hP+C18FEAeRPhb+ij
Sp5QxFHl6jz8gonHJLVrHxRwUwxPETOpz46dqEp0w37cd/hHpXku/i+i/m9fwtyJzPnRJRqn943Q
zlvTuNOlmm2Iq3XI4CU=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ifpXN6gIG+2a6USQaHVbTjsjk9vDezSrDz8p60VT3cRqBcFX2LD9phk1WcldTENzrj2RJakQZzV8
TDQj1BPGgr6/9w4Hj1mNJBWP2h0l80S2VU9XMVRqlr32O+eReCyj794uOsQDKAuYbQbakxBP8I5d
z4myF5muFsnbvA47r0M=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
cCTbdHyTxz2eygqqIHdE/aqcNN79CGIpVM5WA5WqmhuIutCuWaz38TDGtjlkFWWXICSuYppUVfFM
nURqy7EwOzcON2k2AVrDaBmNgqfkg5bgoZzgqOxAyoPbq0SFKYlj0EsCW+VahXAMXrF2ew6L22Ic
ZtF1V62GubiDzOioG2McuyaoQ9Y3mTb3xnm2uc7ivuBXtbT9+xH35PGDDD0+d399XNLVGA6Ff1nV
dRMV0emrUyRipw6hJ/SnE7VRSET1rymhW/9OvJT0417BUop+Wuq8P/2c/IpHIgFf1GOxk5QGnXs7
+GE2e60a5CtOq55uABer95V6yKPqZuS8FN9EWw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
pGEOC0LQtuy+6aWJy7U50mUhnH2HPXhQZ7ROJ/xjLhwWO5TFjBB2ryrtzDzuixOnQTxPgBMyIwrC
9gq8CrhLLbO1veRdtRJkyRIPfzdFcu5fiNVX97RkD+jmoo7/i/y9P0hJRibNeDbDobQZuopD4jly
zgHH1UEtmLeSb/vD0LH06+f7I+mnAMQjexFCnCRy5wpffn0OqDGcZRjN7LlpulzuN+9ZRuSTi4tb
++8aPt3qBAKWhPdIvLDyCkW6GiTCQo7VVOAOF7xdpWr1EC2mxUZPjN3bCbWHW9HhGdsO57CGkyPb
MAbEAe9f8tsANYv5SAjaUoAjBIZd58LJezS43A==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OyNez7RSP7M0//zF+E54uQV63OsJZlsjDWEXlxi0YbpAdRQ8eaeSMA34F5bpN2y5ALLOHMU8CU+3
G8CLbddLs4pUjJZy7h/4r2ZlgA8ut7wk/qXdmq6ATFpXLohWv8ImY4CvLuLPhLURWPo+IATh7Tfm
myX3ZmOb8ljDji21FIflUYsc32Sr+ZDT0YgJdInSvhNymCxlH2QtMHJYnLOYLwYvlckwa99KuEMw
ilsHYPCcdRO+dNarj7J2zdAO1Cw4uIL6QZz24liNtXxdV7oBigY2aQ1mKuyk8YIoHjmKki3Glrdl
RnnWGdoPIaXnFlMxY6gkpWKFLuOlPJHZjvUrBg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 151824)
`pragma protect data_block
f4KYv7qMCu4pAJNp9gzRAL8FNtUOYYa2c9o0aNNKmOZKo65symw2HiKJRbFVioG0vzJzilzFL3Oq
tui+ttpj9wkDg9WuR7kWOSi4JZZi9+tq5kkOjX2bLlTkkB/NP7p7UEgn3bX20DI9gXx9ga24ZSYq
Hk7881blL1UtyBX3xh0pFI3VfbY0YLq3spkeJl4Eup+QhWBEKkWy8dXTEdRqsWNHqULUhRFVDZKx
DKINIwtCywaiHTnZjX6vKlqpLIx8w45sTkmQTzK7ji0n7FbraGDASl3zhyrd5LOMhhQXKG1OIX+6
O9CkDCiyICLazefjb+GYccZg9wYKDQTgWeV7f3akxIcxbR3/iRHn8sbd83yF+FyVtgkoSOyVuLgt
EFn5qpxM8/4mmem5t0LHdMi7J1ar9Vt6EfSAjRSSo2wFfubv4Y258uIPTdp1NnqHyIT7dZ2xbfIo
Rbxz6e7U3551Xj/AWpeKOWepEABrFEygHpnYbB+wWW90XZes5Py1cLtb7G9hbWLhiL6ZAbFAtrAM
MWWtkEbappJZiJ4S6/kbu9ahS8E8huTpCGJSCHWDnAaFYXOh10YCP2fM19JLzXeCnJLkeChpwQYk
BJw5Exp8YGLsDNtxvYqbIol9/TAaegNqpuL3kf75ZOGN9/aqFjM48LKxr48HTXqlnmC7KoUrghF6
2XMVkwFmvIYJvwf1fUoqji9YIscAUKxFFPuqGV4MSslwIhUgL209V+qlPveISjAbkuHs4wY4Oza9
RA8aK+Iw6ExCn7CHEJUAMSBgGkF90smW1jf1ndqpkPVzBtiaLw2drGovM56k8tnUIbxSVp0LqYKJ
LB0rncFIfxaAxNBMf7X4a7CbP+1uTKTR/FMdMw00gITbrzoG3o3L1zw55c6eJfvvL1tQmRaLeLr6
EEFVXtgRNxpuMvefOdCXIpTLNc9ICMxHmoIOBN/bdSgTkbXJyrWRyzv+651kVLAzrhvZfTtvnQUs
jwAMPzu06eWy26V8cuSu42Opc+4efQ36kckcAUaS1kwGKoE77Z4dgSoM8jQmFRDuevviC3A4/eJ5
OcaLj50RvOhd19Rd7ft3BMFsp4SD33vbjcum7U8hKBzm0VImzKOONSj2m6MhlfIgb4IBPGlgeXIU
FCrTGjzcBDzAtwxF7PzLjCKQgd2Z6kHU9Vi91hk9G5c/BYecjjYzgzdLMjy36w1wbue+wiCukUud
pCb6hppiU+XqJiUC6E+I0GOWBV2GYTb18N9R7MunVQCFGqs6EuGvT5Pfgp1WLB/muQvF6edmkeh6
rniPMEjqFp1TroZravdMwgSbtPLFHaJChF5ICNQynnbmvaMpmHt3zbR2NJw6sGD1ybttt4yRAlmr
52AQjYRMFfU0PNUb3bE0j/ZY7yrXAMXaBncZ4ZqTwcjFQFJnKsLe79+5iz+L3HcEWtjy4O7JOyjV
2ZsK8Kbef31JOZpKY97dYWIT8lNLZlY0Zlf44qciT/IvWAscwnydbNP0ThkPsECFHNR0hJJjb/SF
8hJcZXZ2iUhDBrD0xHtLRzy9t86w6lKEJNcgKny6jo2Qg3kyYS01wrOmgB+W5J1FatTx73nqIuvk
VZKveMhXPCXS8Cu0bws/tpXnNjgcCrDhSC8FAx6OK0LMgCJ4w3FuKGzFwclciPhRWIbd6CUExBZZ
Im3wfRelAxL1mdcblrmrEydfHfjKOUzJI3frJtdmv2wCxZxNYXmbg00JEOM/RgMpx0rTVa0HGf/6
RU66ZJbwiZFioGbzEA6uC7RNsZAK+gpeOncuChMpM/SEZOsdVYQ3tr5mm5H8oepaS+ywWXFcGVmO
2o635Vt5XB6iZ2DAS1LV4CBMQwoj+Q47GL8UYI7dWIFJMbdMvps1xKw3uW6Fz6KwIR5QSIDQ9/Oy
FQ4r+i9DKrBmS8Jro9YpRbTNNfM8ckusFmUnb5I/Fl4AymrTXv9ghDWoMr0AavPG8LExUxuR5WWi
IC6MEmmlLHVAo9DRFkNkNrVKSaGbiFoRdAqq8hS/ElzrgPQqWwPPbhizfz+MWa2A73os+2YoNZYO
xjKxbw9vHXVJS5jjqFlss13siECCI4juk5/uOkw2Wtw4v6PhAe5wI4VOJEbnewCTNvdR7hP694ld
j63yyJGcPqamAoE/F9pUS/qHy9rZ7jrHZaehKQkSsmx14CMI8hdvQ+pBeHj7GMN1lvv/2iVI57p/
P8jaJlO8HHAyDMBHPnf6gGb61TCwENoLEOnRIg8L1YAdAVfhrTIeLfhjv27WFxxNDNFgzDeVnep+
5CqcCNyLnDlmAS9dv/mk2+XYKGm5ssGZmllEgm5ed5MlFoTAZua7J8fLqiKiiPbfad5NhEzZdBXj
0VD2XSXbj3Ly4z96yyKfcbjrQPqtVtnUrScM6JdTHlL4bHduBP5Lqh1Nw5CEUbY8apaAohMhU0cy
zfKX6JavNQXZECX+gKDJW5y+nl0TEcqUK5d5TcyEj4FthAQX556JobIv79QvPXYgklDxNzRd61fa
00sTvfinaqA+i+D9q7UCKnA4DaNXSi1nwiSxxWzjrFUxAe2UMMAo7Y5cZHG/8/theGQdzmn97Zk+
wVunmfw60KB/dqPePjxS7JGOQlAeie+s5dEBnIsRESgdOkkQ5BYWWLzmiOMwC4qOuCiT/H7QeDHA
Z2WdDwr9hwL4QDOeDj/1ullW1/PMazQL/EG+gD9y+0dwg9odK0QiWgnkpctVCoclSmxhJLF3Uza/
3iLqUGuKHB7jZaHdx4AreUOc4CzpkJT7j+t3j8A+dSzsTIXOJLITmM9yTLNkQsWXVLs9UnMsRL30
QHmMLtSMTjjYeSDFMk8w5S8GNhYmh7aWh2KPLF4SPaXg41G+KGVcdyJ8ki6/rm1VO86STWzR9OWT
HxuH/5513lOCQSPovAoo/jwAI1kk6DXy49T8BkTf/KX/MdbxCitwU/Pmzzj4DBVUdmGuvyJoBFw3
Qx4HuC5KNLmq78bz2zEiOB0RV/DQsFkCHqiRc5BChh71dQSe5QJCG9WJqgS5luwVS1eF4zt4deQ2
9PveE3WlLFTU5PHB2zkOhVRC2yrHLyyJESWMeidwedPgtbXGSz4cn9CD1oTrdw/vjGs9/qvEUtp2
+ZPyYBTR+gaz8fKm8vvIrGoFbUQzB7gv7NC5M26YDYWYnVJNFaHFLlNWovlKjOKbLjE7hdiG7Jj2
q4PmmzldLF4yVmDJh4s7Kl6+BHSqPs1qj9e69IicvwD2datyjFxJ/cLF4PRixrjZwSgwdDWefxrY
6t7M4yzHBQpbuKxGbexwe8ecKKNvxjMvIxG6xCw/Lz8DN1bf2g61jfHYoMyy5W3PQiYPVZq4NxjV
kn3CBaHNrSxfStYwFlzXafb3A/Ze+Z55ynU93CI1U4QD+gvEHZ+fREok7H6I4bWepWT2rvEx3dZW
/Iw2dwlb1WRRpXpin90p+Qn4LSOKIcz9jE1m8hQRAPGx8Kzu3G6Aa554FuUrR4rHPmY2OoT6OAvR
RkTS2bW2W2CPCUlabyh7RtniWY2DRi0s24EK7iEJK2Z4Y4W1Qz+PDxjiZehAFBo0fcUJb2WC4VKC
reNFz6I4iRmt5w9bWh8U4DSCl/G/99EVIbHjlQcfWe+C3oDrJtv8C3waInsq2OuWHKCtWXzpps9Z
MV4q+cc5QPYBrQqsUk4Uc99eJzNTnW04Q5pmoYv9lpsLVZndMJVo6DvQXvdFh6pafWFXri6aKxFJ
Hlr3/vW11RZbAPjQFEjprR9tnZVZydoM7wEJ+sfbpLugtAqIpIUDhQgyWRHOckTRsA3FQBV4hejE
TvAE6T7Du9qJDA0utun16g7MaxobCSJClecE/1YnDUYMkvXScLt+QkSmCr93jqkah97w1zmYpcmx
D/aM6Kgvj2jHtwSuQZnvWBtyPxvOv3ozQrFyIlxJlQIUOGy58QwBB6IKkMGLJhZoiyu2c3y4TYky
ys1mEKYaznD4sKRhF0vAVgFYrVDeEw4V7NxiBYY8T307agr4Cpjr8eqlTOQXILpkl+tUzPia5bAD
Yo0B7jgxwlVHCnfelpMtpOjCsAe/3lft5JkRhu0ggZJb6l1k9JwNK2xAMTiPBwTVoPH421lC4GrD
obAXwNJmhn4X2TSD3VMz8nyn5ahweaXHIV0Io+j0WB9teeMZVnSM56E4X8lwcv6oicgLN7FwP7w+
lfaN32ZTX0gYMe22nVuVD0v6jBlh/lYq9Mv6wKpzW3bHJrdZV+DE4omZ9uxAzHzP/7L8kQEqak5r
I0LGoPz6H2xzY/ssIWWzvoZnRobpxySKi21RPFwDN1mzPdGI3MibmXGt7ohbVDa/8UKyDMCdTVcG
6fkg6sU/EPplSdDCYSc61nj4ucEglwRDM8osnvtIvfsgADPM8OZbXs3NS38iuJQYmsBvBQ7F8pJB
k0Oaa4GHyscvjpLVMx0vJnhwMh/n/ijVy4WbEqapics9VmhaNZIoI8VrgUpmHT+NOXG7GPBaebBO
PnjDZEEm0W1XcCXqwwUniBZFKJQgJAbF/pYNLaTyPVg+35jSMkJkV8OFfCCLk1zrPUtxZni8mXU8
FNjsiMVUaLAxb2h2Itnz/SyvEHCLYpUjNb65U2qp6fygj2gLNzELGtqLqd1o8Ak8vOv5K8AaoDZn
K4O9MQjlo/avTslSz+UeqdslTHxGtLAJ35faX3fYtjZyNXgV4l6aPQnZSjYXQBLCQE3zzdWfA4I1
OMAYim1f+1uSwySNBAzAPDw8D12c429ekSBu83ZMPikwxBkZW/Jb0pXEtsGC/iV5hqNpPIsRpf1J
/tv4yrCCghyyYIjJouvTCuIfuWewC54F1iwP98IFEyQe+x9pkhGT/KYDcfnEpdxRat0nCRyObV/B
OXhdeGKMvazdP0ZNLHQfduNe4D+ZUSEgo+acfH0BPqUsAsoHpds+/P7uNHgUYWVJDkcbGmMwIQoA
skU7U1d0HG3di/eQ/hfVR7ybWOn/YhItrRs4WpJ0nvZ1Gw33EnJxRGhZCXS2RS25KB2S1EjK9WF2
DDCZkL/KEosFSV+MJt6+LpI3StUQbC2jjM45Xt8IvyEzOXBBHux6EYQFgIViPWZBTk2nIWExYLYe
R6ASOfqi+iXZVcIrB49b7nQqC03gupCHUGZ+K9xiRFKFyumohJ0SAr0X2xhuz8rMqzGEpgpaLjix
hNWusIklrX92IW66F5EZIJLG4ECf4rV9eFiPYPN1pNBWO3Sr+u1Phc6MxLOHfQj8foCGyR+TNcfS
Xp2lkvF+c8e/bVvdlVLZfmZZIQrJjM3Yk45OfSkSB4nX7W49llk/KQ5ICh4M2OCLq6ayit1k3Uyy
t57qpzu2N2dEnoHWBdGvWdb+Xnu/rrxoYZ6wXV97lO+Lru/cSRbtMLTH84z/DteB6x+68GNcQvQc
zqaHcSt6OtKH2uNdMLssvvg+7NyYNVCa6vv82VkuHIlMj7ewpfl1smokRu+TaoZglawFYUb9hPGR
eOgwb8lvgUmoijB6+VNe/WHzfJirc1o0wdGsexTH3yrUa6GWQ8O2cyCMxsrC0v51cDhrDqVXOu5s
b64YfiRX8z6OtiFwApWvRWo9Eue7VYsMM9dXWxZ05Qxlt8EcIvAxjbnpusuhFuj+xaGYIl+Jv094
0E+3NguKDzXJeu5Oq+eeLOl6IXgKMKtilZXBpvSxuKHBpKi0MTMKg5StcoOQPv1nL4HRrhXd5XoL
gjsa8gapMbV+Uz6Qa9C125/9KlXkB5RYNH4x4n4RaldKTMkFBdJ6busUGATpPqDgeRssLYbt97fk
zVS2+l5Pk5m1y5D+vYoQQVpX+p8KZRQBNqKht6Qx+LjfcP95c7KgGBAPViKVKAzcu+n70lhk4Bi6
xmIBi1RQw+A/6xk5FVRKdUXCsuNsyJdwcoOUmL5Vpr4UlARdDsuODsrlQ5KIk0+A4v5R+Kn43vOd
QrKmRQnXCSDyDisFX3/MITpGieyEgmEx5HCVAm+RpLtQvgdBNM/wzcw7cEaQHQRdnIRhuOeo0FxB
2NMaybBeUIA8u6J1Vk+K5pt43P8V/kJJYL0/T9W2bhEpbNJ0pAUrLCUETjjGPrO2Vb/WF2TF0K7U
k1Ie/PQqOcdpNzVWn6cp0ptPe9dgVi1FoZeutrxDiahl25M1FKriGBImaX5pJl1tl4/Y/G6J6qQv
y7mcECzy0MQ4FQSIfJq4U5IXXC+ABsmlcKXQNGvE7sJnriMaQK02c3q1MobzM/Rvvf78Id2xaXnT
eW2kvKtUpRPDS66pBjP88C3t+LTEde3eA4LA181vsISlsMtXZjF+DHs19FeMpxjssq78A1riMgU3
LfgVATFnUuQ2WIBY3SkKBecKBN02PB5VH0w53gfr6QASpKW9tKcPMC21N9WEGfVeVUl73r9/JYZX
o4Aq0mKOca970yxWySINmJE8iMrGaT7Sij+sRC/t7hMJuHSiLcuD8JFKOXtYcT2D5huZJs4tAYbN
Wur+uNrkeQxF4ovZ+vo6XEYE5vBoCjzUwIgHduI9vqdcWHFoSN/kaYcEyvBO5gHEdikB6Ff08mWL
JQJe+oFGJQwVhOll9IIvIeHiutHueE/hjoOTovlM3rcqlwCrECTrWhWyruf9P0wJk7nKFmBB0rAx
1nVTb8pDiJRwEXoBio2V6TtyjxkdvRL+IBHWmUHkXAczHDXhvztbqiUGgWpaTgJltSry4f60dGH/
abC8JZr8Y3ml/ynHnnZybW7ktV5VhsME94pqdEY0BLR1egEPXVbXlRsO3GTsv1haJixH/VyvdLgQ
42tjuDmnYg80T/luRTNfiM5vhAe9Aro+jIeg9Gx45lAUSdZ+Y7in/4ppi1agww6TeUP59pcg2aFj
uQAxi8dRXoh+E/7C+llNwx37sgHSDLzSz5WvhPEQga2IaUX1je+sPb+xU+9KYMro4IeLFwHRqNLM
OG14wvvgrP5FeXZY+v76WAnsXt/wMGk8GLo2xaawTYxUZLAJF2RIxWGzLbI5R6mVrZuTwcqO8s/+
xE9KZ3Js3SLjyWnztutIzytGbQYOGEiDz5c2fEg6hNEsSIyKPH3QHKrGuvVmb5a2b+/U1v57uopl
NX0Yx/ImiSWtDibisuydm3y9Wv4sddvKpBZ1mBlE2zqGcWsU6ZXVDAyODR+N+QNBuhkDISAsD4bp
GDGf9SD73ZXDF1AXkRvp0JVW7UXNgC1QjnVHtDLRNu6UrKYZQjoFkx+kvC+hVZMYOP4ZUkOqxMPe
JUFP7k6yrocYhgI/BJslb7OvWISPRP+gb0kXAnZGxhCbISIqX3IES78OWsyGFlFtpzMEGCejNsok
dOqQsR9bJXbSp/xXIyUPB77uU7DvQ46ECpjMmgUhByMchRYNv7lWL8fbcgpZo1780jzqogKsB1M3
mPxFJZSdJvpBmfm7SPGSZpNWXX1/UvquHITbdh0CM2FR3lpIYnlnK7erdCGB1iiXGBYfzUqb0aL2
aKThFutOhYZNJhFYnu7LrCdNTdaqz+br75uMKV+O2ksC75EHG9ZU5bLRDvPnumW9oj0Fkn4e5PFj
5neR0IRuU4u41L4H18WioHC25hQQKCYXbmzFJbG/evk9rr7MfnwnxuceoSpRKhlhADqYgoY8HXIP
BUqxKNnGneTlwORl5FoAQIuBB2i8sCRXU5KD8wFOwQoMsyBwcd5U7hPp0qFBH7IZIgT6G3/1Wtn6
a9R2q+DSngmdzy3reRBgReKiDyqC+PdqLIiUhUoq/5DHqJJ1b0DaiiS72dEF+YYGoUWgjmpS1PCe
P+Q2QYCVhfi6Iiwrh8A1hXuQRyUCe/ejohD//DpRjdxSInMivDhLUYXqoiVurdCBq+PbnwjAP3Yl
XRqBjApR3ac4Xya066NFVzdY1gz3Xy3LJjcqToBrr6u2M2+t71+gPOa05mEI9E/37VyVtNQNl3ew
VEyrEC2yIbRh4zkIz0ERelqMW68l88XZNCC9CJGbq6I4xvIswNKAkokWR/flFpXoW2Uea+cLGkmL
DKA6CYJWr0RbOWIZocvPX6E/rnE4d3vnp+axvG9xTNiyd1GpYJgEztrBtJHJHjE8lDp+u+v3ZWLv
OhI7oPexbuzdtuar6c+m3arpe77dveVPvGtpTp8vz1BgjhdjK2+ipg3gbP5lgAxHC1SvkHkFfWHD
WlA6MLSVVDRBZpUYr4O0gt4pQoHHXN8S3INF4ypeaP700J/HQMcAGCcjEZQ+bkHo3dX/MuFe1gm/
P9QG51pLWUrxuaLSV7BW513guaxM6iRBJ/Y0GgWlfBfq9KqVsEKLZkq45C9q4b9OoklVg/GLoolf
V5xfUw2vI6q4zFudRpvM6owbAU4NKbvfNPbBY6I1ydJ7cKvtLUWf1We9652oc7RfwmDv9MEM2vS8
kQ0xKdrXWsJr6dWOv1sVEnKiOE+2HLWvgJfbJ/vE8X/1UvVj1GEjpqHVHgJGmLuFRBw3D6e0Pv3c
Dryl1q0Riz+zavjaNl0QQ1dtX3ziQHjby8EddKohSx2Ht5kj/lkeCRz/VNgW1zb8q0DWLRM4GAEZ
aEYKIYVehM6/qoiQioKP4qocpy4gmycVOaOnD0QVD0X19cfepjPs8406ngAUK/ak4/OzZHv5tgOo
qiXjXk6RxaqKRv/YyL9pu1WqgcmGXqANOMHgmdKCfj3kKIlbUZTXbEBt+CGmToxpSohAMd0Gqz5Z
umx4p6SMCJkLNgLMk+Tw1U1D2IsgyRHKp2zG103xNdFOsVCVpJQzm1sLmr4XjdXEERXYKnAcXzxS
SpGVWpvCe1Ol7OIgK79XGHjgWgsYBnHvduhdORbE8pD/7REqFuJkqwaEyQMsIUpDk8fjO+QhgYOs
sYn3vCHlva3CsVDRSZHGvdNcoCd/eooMAhfVbXyPylb0BQdpaVXxUFPK65YiXUCOzu/BYorjZnUE
F8TdHixBO07k8w2vbde4IDnDZVieUMeVsfxs5YiaV3Zw2ZD5Y3Z0m3tg7upai9wtmvbNjOXhUNy+
CX8Jycr4BsWF/F9xCSYNoijFnO08UElFGnSa4jnF0RGuQLzu1F0qZCwiIoomDccOyeBL6ThEXJGO
kUFi086WlpT0Xn3KRQtc3mEOR4c+wOBo9eJMsYGtdNbSYEZV329nI8t78yorVW+3hr4aaxoAtWSx
whX9efLfK82pwnOiordT9m4o1G2zXTG4gZNG1YxU3pOaLGoGlJedVd1UKvZ0n94CVMS2JvhIFGQ9
fRKGuUl39l60cgbDc4rsIFdRlaUVuqyRM9sXxo80fMmcv1Vc1jbmochU7madw7tmilKk7qFPiFWC
BYprzOr44uXK6P/dznSoPAVRcJomdF9UJynwl5y/oO+c64nZL5sEToJ3UalnEnIdV5veiLbz8rLh
lgyqr3+N9CpmrofgRT/Oo36jePWnquf4d4qlPlBGugIik/y1U54eKdvAf8mZSMKkRnhFEnRIqRCo
tgBvX6LSStsJ1gmFLojTTMLKSfoVY3JFzYmxxBd56TzGQ4uNq/l/qmYaD8FWNy8gjMrsot+497tW
a5VZTcOwtnrTLtNycjYyRhZr5MXmn2dNSJhSBgvQmm1Ygk9QA3NNUSyfGNDP02bD5xZC5Scsi53s
neuy/nARGywpv/v5o5z4mUwx4MTYK0sSOwUxkW12SjVPavwhlTaDthGBixgxgUV2frAaAttyrv1Y
BxxnIAj7JBFfK4u6tmQQn+SGpxlGR/xq2O5yAjZIYscYsJ65A3bj/XPbPQabZ3kQba/vDfChvNw4
T7CJx3zq8MD9Ols+pK9FW/ALDiMgaZv9RRWsF3Da2UfhJTiqm7okRZMN0cexGBOHcZV0vIGwBrDW
G1KIO+bqxD8Zz/UWdDeJmhVGNLP6vcj26cdkCh9AgcgyDv4cP7xpTHz6x3TZKbs8jq417rR/LJ9y
cYWG6k1tzqRKXMIDzxNzjt2yLDMkGbq/V5481x6VPTML2W82NTcHL4bi+ZQ8psxBzsbKcuC3Mrcb
Kl8MtzzlWnxyR093Y+CAxz6Y0mRsmqnE6sRx8Cs0bqPijlSW34P/Mz3qRb9U7V1gb7xDr+8l+YLz
4QxZnCZhDuvVzT4eFizOGFcjX2cVoHBLaznlHnR1vKmurq/H+RyhJyh1ToYOwMYnrR65IQO6R2QS
IUKfTbEyi/0BIaY/FWSevYB9Gsyu1IYlPS2NtePDY00Na83BP6MdFp/7NBo1ZREDOluit0NH+MmK
RwXOOunhahlzvEOPkNZao3noUFWTYC9OqFS+DWvrTZE0D1HT2wjKcKnv8JwDkrgPTptkn+HvFEil
k1cZiVWxELNaAorspfxNeTsNR5czuWfsdwkc6u0Y8swK4Q3wmIfB6/FcXoffmh7lfPr2HRX9rgUT
EUD8DFtsjir5XMhQ1mLJiuK5R3b6yTEdkyW4REhR9AOQDRSkECrJaylAqAsxgHkZo0GjYSUWBtv7
zokJ2lQgy554+VwkG6sKT13AXCKJzX2S+v0gTuYOuRLX4HLKkEShJa0LxYI+1P3EYUIAtBcJpXjk
g4/YiLONCnZAmyiCm/FcwwPb9XkavVtOeG1+GECqBNemkXhpghyD90t1b/Zs95nX2kKhfv6pAxZD
Gr8W1pS5dc6VhQ4LwYTC235wNO12v2TVuV4Rk5SNPPSWyBN/toa50R6z5GVp7g5PF7AHfZIh4qN4
ysaWIOpjqNiYKJuUngcpWIfGv9ldZ2hRVmZN7eOijCKr22DumEG4HoHQyi6B3K4qZt261BHB1iQ9
UIw/oAx9WxkvQKkci9PTqKlksvlOypTRoXq3BWL86TdEjuu1xToYWgG+mtTJdg9LGGFjnhtF0DCm
8JN/C+XAVf1UyHOxlFznVu7zsG2elrHWwYkgjQhy4XbNalHKBgIv6oJlMemW6rK7vrv8iUPbJ8MX
AvGIKGNpy9W2WAqRwrCczSw6a0imiRR5W3Iw62VtMESIDcuT0UHZQ/eP59oKmtGOBlf25C49/3KA
991g3dXx1K3nCNKeM3yEXv2tWw6ZLeidZoFK0xoTMUkArm50qIiajNHnlGMwerZsEH9TBPoVKHbF
goN0GO/gpua4/V1OpPCZT6LCwfGDytBuWInoSh0Q4gHaIQMNOiG281kfpSm4Ejz+47qukoTlyl5G
5jaQLQggsw8Nd/F6ARTOFeELqh/KXH5iAi62IlMjrSrtGMwlIBEHVij9gXS8aC8uAMZtrHMqgyKy
nwL8tazgkyKYDnIhxCgXaNeiAu1oG1FldJHkQ/yE9VrfqW+IZwcoiqMzfkCaMtSqylEZxcpETj42
Df3Q3KKty+eaLc0U9CQOVgKeefoRP6q89hHBIV1byX4FApuHYg1bsXBCIygSIcZ7+WhdkJzeqF32
dz513Kqhct9fbTNCq9Y+VrvJqo2fMJ1ji+vaAx93QG3/io2TE6qsqf7sHqISwT3XJwq5WJR6+0Ry
Z3fFkLxefPUnkMrisPlt82tIeYG9iQjtaGvlNfwf/aH3mwGMwAgS3Hq3IRic0lNyRwMwC/Y4F5kN
cQTjP9slfDU30k7Z+HQQi5UxYsYx8gf4Qkm5q5Vj3+kALVmOgrcnVk3RWH1Oy4cnBE8CLAaeyO5K
CTOSENGq8rxbnkCVhHkfaTGp8s7neEY4z613RtICgElXVUoGG3Oky/xA/Q+PvWtDF+OV6PCNEyN2
fsJlI/NmV3rToPcqC7lnvNDx7WPbocKTdmgmRG+ULQ9m3EHHgeytZ2+O4WvmzUEBuI6oFJt1qz+T
1DZQfu26jYWWW6GNmBudaLK8JON6kKLlBHTFqfbtoTvpofhj2LZxLJYNOUN1RclWo2dPSHf1I6I0
4RDn3pmGdj4hmoqBVrfaeIKPWvGfLrhQZUOhHj4lx9GackgPt32BbIgQbX5+6AUlrwd+wk5tFOzK
z8g2EVjdkbYWuCP0lYhK5HtXcm9ffLL5w1hvZ6l1NdjdIms86dJ9iebbKeeNEbwUSWcHnQlbHSvy
zd6SEhRXuLuOwB/6JXNRM/ROlkwKNNO4SKmASWH2nIcdz/AqLv0pFpQ6Ozzs9kHoiCrYqqnRHJqS
6/F0CT2JjwjlcRZSQsBJttMKxCxPP3iIGdyeASDXhk35l4FvYPgN5VOWu8R94AsCol6RuqePFils
aatRwLRe/I2Fq4ofHsmo7NWDiRTqqlBc8VCKjT+5ahmjXRSODA1a7Q8ojm10hq1LSNE8K2LKM0HB
Pv1mhgGHaNNfXVYJnOqhuiADsNvkSAVs7lSS13kkz8d0U/SJ9PI2ZOjENGJ7ai0YJnFK6B5adwCk
CVHCwhUpTtYMniJH5YY1t31P1A62r60vRokqb14+UA7z9xGpntGhyLkDO77wK8glJoU8/BhC7NGc
s98NvGzlrzGS1vETM62pO/LGM2WHM7LoQrM2+vgzN+8I1Tfmj/JGfu3Y3Ad9RLnwE9Ye9eyvoCXo
YTD/ocdsyDYTqCtUuXuQHk8HxtPImfk/PcvhTZC6e51vQSxSoRpMepECPhzjXQTieRFrfxFt+GDJ
tAcdtkV3rbMQuTJ1El80W729Q4f9poE7fti8/o+7D0yC/EQMDNrCyagjEFgsiIn8zvv6SrOPDDoz
oHMIQIHK98NJAhG2JIuv/utrRsUHRKQ77IMOhltvqSKvPN69ZpCvD/RzPIfk4BlF5jHwSvcI3p+r
09YM73QBEgpMjMrC4/ttYXCxfW+4MgEgDjVv7t5TlgHVmUA4S9bKwwqz6cVqJrhpcz89OaMB5dAj
nthN51q/yNAnMZ7u6cMrpRSPrSWwjrSSl+vGxJP8J6V+cb8xy9aIDp2hT3g7VgR1Y70r6u7qWlfC
o2TqTTEMKd6PjWm6JKUWh/fJDpuFcGdGcHydrh1SfzZpUhQqwr0aLKZ8ORlcMUXIubKTqYNW8iLp
dWeQnD3/nLH0VagH6q7/xwK/GWr2kbI6/JqkuXL/vD36mqGxqF2dkh4kbNLOXb8vsdKEAprTamuk
r/HgsnmRjfN+f1pCIIoEZ332RUvpXOz2ul+9UUwRKZVoUR/c56muyuv6hftI+m8f6mNJg0Ihnftq
1Y1QhAdhNyiBYD1wfvPZo9KCu5B+0FtlFg09jwHI00CXydwhW8sMvJhydmNkQbI/C7n4+qjfhKCH
GXPwdmhxhNd/7LiO+qqH/PzUzO3KHsmObLmR1aKIhyRSjSTDh6Y+V0yPdb2jJulZJl+zi3MAQG53
yfZorcqNyj28z4aXJCTHHduWPUYsTx/t/9nTF+5AArQqFVOMimXo1IDo174Jdtn5W1R7Usa/J3gt
/3/VBHNCgeVRpVGAAHVGsIoCNDlhBcfAOxZ/XoExUQjcjoLR2ogTR0zk5FT0RYattDjLDpq2Ytii
6+tV1fIJhexmYbsf9jwowM1pdHuv9Z+9Stw/+z09C+SGH9zErJGDabBBC7/PdmJaGehIOWYxfyyd
NrwVN8+evCr11HPAHZGSp8w3W5JSuEyG0xsS4z4qYP3FPoThk9OK+xLpJXO2NmeaxLTqZ03Ehoci
BHHt6tN0Smsd+sYsf42AeqZ5QXK9XCa//sXPPIpHCzIRXeq7ADTbvvbWblKgLbAi7dm3mBipidQf
J2oDlmazVB4tEnFFrNjiDCpj85XLwdhe5G/Ko+wUZLypWdOBw6zyaPxo59V8jU9md1zF2oQHCSMA
zoJltuIxdJDh6U32+e2CT61hBOj4atWyIwHWXZfyHRkLTFY+YYGHu4sYKoi6mHTQ0vxS9XhC2hfq
Kmstq1P94b2UHkxktideQDbk6dLnlwCBMDETjAcjTFO0phTZw1HXUqeMJciRx67LT1VIxZw2msOj
pqcEBqx2MIKJRN5A/8S0W/lbv2vFAPnEkRqVogESTXcGoI/wI7Munli4PZPEticZnFI/B0KXoqUT
/aFc8IxUubW2ytgdp/nD6ppsMctNIzBQVk6UWnXlO97vDvkWjDbxlt+fTvUFg5hzoV8zXGWy285l
eQkC4ool8a01DEjWj2+Rs/4YPpBLf+W6X9fWXQsiuYahovnKwFAEHH3w3XIs9Q7rAc3P5P1LDNHo
NGA1faNqrRehyy+9GvCGy3K4nh+5tOCr+Up6MaiUa0f/kykf0oBY6EGW5WIU5ICTcUaRjgfwjF3J
9NN08QTRtKL1uE11S6yq9x9vwxX+dNEzkIayfobu6FRcQWLFqSZ9csqO6jwL+valcSWrgllMoXxN
eUBVboy069O0v5rEMfmOI8G8HRY1LYbUqolxk+O1IkVaI6PUg0PPa7sH6zY/+ZwWy9yDlDSamv4R
agpl1gsroo66aWlSHKw70hOOjxNIC/bh8Ylrjl1XKrPkkcpYNq2gh+RkQxvokw9Vp/xK4ZU5DOgJ
2/Lp7HgVxgkKxjlpWLXv0WU3TlcwBLIa9zNwNKFbQ50i1YQ5jiZIZCmCzCm1v9OH3+r+BEkE7Fdv
QZT6/CHDj80aChX45h42fntEl93Rqwu+fgwwT30FgLhOGnkd9+qhkriZmQlmoo3A+/9XPzYA1IEJ
6njhipwy+GopAqNtKxkeh2bOhP+TSZxlr56djrGDbZZlV9IR4Lf70ab9waQTvqEUHeDLAIauVUpi
rSfiJ43n6ThkZ3Kw2XvlLV+RBtVYuJUrgp42RtuKMegVVjAMvI3wR7nyM6iqOghdtz8XtVSAQtSf
lI1lXjnD2VmZ4D+OXAYzltqvvIkAKxlgFhXw6eqPQkmT41VeBPv5sQbYxoSp/pIocCW7Jc7bGmr8
de4gxWNGoD4A8/RJHF6qmbMz8Oco6lGOVJIAug91PN8GdvfbVS1CHOrYv2PzBDnEZn5hS7N8rItJ
3CrQRXkS+3RiGDJVAmZi3sQCeGRpy8W5y/oOrox2erNMjlx8djQAoqCSjaBNZocq0ennuq8sayTt
MvsF4OlnqKTzDFhjS7svFI+2VIT/QAW1cGEiUvZdy2gvkPh25Hej/TdosqZT8AWUD9dppAN97Jav
+ytHlcmRVbmgXxOkCIiWuxb4neczH3Ca8be97AezDWQYsVR/xb9EHw/3qiuonLaPO+UpWHZb+oj0
0eU6cr+gMIShsUMxushMo55kxIGE7pW1JELsHnJ8RkKydMYf7yJtw73PhLN1hgzbUQTfuKVzgxWs
sV4SgFUItCnd9mdJnJxMCokwU4EoHI+v+0L+37zG2uNWGB/6rQ89R1JO/jtTg+hxyLgiN7Tq1bat
7hdcC5q/hz32j21a3HwXBDC7kbFnU8QZVtWoj72sl87OAlVVRviyRYC2ic8+vzg5fKMP6TGlU2Wt
DplKMnXNiCM+2I0itzHj5y5RMx9cX0jKjnInnL0uvZJBCpzQAu8l8KhL1f8IuBipCQMUPUYw8Fw/
ePZPKM+TB5s00Kz6nGepPzRqRn5/7YNEezAfLAub6VaUBVegPxEs9h2uKjUzTdVSqVwY33rZc8fB
UOTQCWz/BUPtHFwtiRA75KReAYwH2az4Ka34nwNwtCl5vizQb/H/QMdm59knVsBLLBj7wMoO+Jee
duXcneXV/7T0hCmk5uHCit66K55IUrGojbucInb7QSqPO7FfH53bayJjPKquHYSQT6IE+c7X23zW
M1DA396O7Dgs61NdiCMxITT9HV9rXPf6MajOnvg9BdZTdWXMGjIdD7rwcLPIX2kvgi0U4ie71Y8x
WHkjQdj1JkgsHcuNbx1MH033F9dz/ukb6sWyw7UrTpK5Ps5i1fnlxzXozon1yp5AjK6pkP8ADM5d
HyfS+onVZ+C7UhESYDlkg+iBZGIrZUky8S88sf1d2NiOww6dZk+sCPGur7FDqAt7SKozD7rpRPA4
liibREy/8hbzMNaR2fSsaOxX6dmXgi2bnzbyJCsOva/L/K1uSNn2/8t5wW6jMoqtuVHt6YNWGeUe
1G6aYbslWY7SZ8H+pgKDrWW+hO4fx/eNqOSiTF6HLKlMoHLtOR0QTQE9At2gb1pG8OBcH6Aj9brI
qCj51n1PztAmEvyOx81csQwuopN2jwAOIbhAJpAHLZjhNzw24Hf0H4pc1RnkY9V87V/4d7DUfxzB
ghnQAOEdpKD/BOVTCnwBdXriMeyElvymiLJFJ0+9PBCr0eQhepsDoynwY32WkijahDonit4OBQx8
JANVUywepk8t0zJpCC3Dhhl7KE2Rc+fI+GUR9ZnuhtV076pkRKUT0ezmDG49Er2uGLq4AWaDNmVF
tR0GUCYrWaPqjmNshjV9tEsPUdPcCNZ2/t1t1N3NEzPAg3HiI5khmQOM2txxH7GPlpXX6y/2rgZM
rP6g+UFVCoBipXz9LG5iGOwfBCqRjlJVh85m6bLzXTmF30y/woZt1jWO+TDguvgaylrtEIZiyRPE
y3Vxxw3REFph8GtyWTD2EPx3SNMibAR4DWh3ryTtdYkfHuSMwimnDWYtKVFDPLqSKIiyeKRo4C+w
46ATiGZ58teFrTAgehXqEIvUc963wtfCPYqYvwW64Bhbx0/aenMXA11+TCJ+/BjFVVsurVT2b4/h
5kLBRAN3ijvwVx0NBazpeL5y3Jk6Xg9CY6g7qGQCQp1aHJDrdYib1NtQkn4vcKeQRZ4y5eNJ6nTX
ZbUvGrilzmEc0Z+8Zc9kAY76ylEodHGFsgdeyo906JewnDxWRQrWpOTpf7gq2cWjHuawNqrDybbN
CZorSRhxa3q4pMYl/xkaHt0X+beJVWp4xl414nRdMk3negjDVFAL83JBv4jaiXZZwdfYfZhYlycX
+5g0LysRSejDtvN2z/3slWJ0WNrw6e0eyua2l1+oAbULWLTmVoBc6MfPL++qGXAORonIcwfZneEC
pwDyYj/FP0G09iqP/wDZz7aU0g5blYYWJG1NK88eaZXuLqCcBEI3l7lWaiT+2ZpgfUUjjrEyKYzz
LAKsvy8q9Zi9Z6GTzoq6Id5JiNpThuibFlpxMEIXmHHaCKzINtPXF5So0R36Kcb+REBOgp7A1f2Y
PCll4U1SiCdrq2c1w8VaEGpfGm4vjE2kYYQNeGKyvhTQy0ywa6cqwRl1il9l3eiczxxadKZUsdeN
mrMod1VhxH+6syi7MXpiIdbN+49hdKRJHgpkyEUSEPKnMt7ed0Q6CbyL0TkNZQHNpDPKd0LAcV1T
IfVxaVtQsmlyppnndWImVzm6jUTz2i2SLrKS7X1bsnA5NNHCovls6bt8yYzg8ZsgLCR7aYKxmfaN
bZNZGu24FkjxrdpP511tkGrvdjrLZtrv3P5k5cAUOwZ7Ti1R58f5CFtrxno4Nl2VouCnDnVFrEAV
2ujMgTpALzyQagjQ+woTXwmaTXVxTcghYGSFsrq+tgaOvxT+UHskjf43FMV+qIi4X1X3OVLlXovJ
P8pl+m/VCWkW2SxMOUkPBOC4pumH07B6n2m3ceADMXLeWJXqbGUdj3fhza3+2mAsBh1sRd6ZpSp8
npaXoMceiwPC++6khS5+03diaLYgp7YCDE6bVYXhmOxn8maNHRGraaZKi/2d7SYublOrlJ8vyYcr
Uksgzj0QsipBxjqdhpbCqAr1mybeYe/IZN3Xoo95wG394bhe1MLNgvJEjKmOPIgLNW6XyE/OiQ1r
Z8FRymMh7k7d1hQOQnAYr2Zdr7a4j+aJGsJ5b7qe6ZxSqifH/b3uU6xVFSNuYYr01PorXDNnjniK
HAeODlv6uKtBiHpviAsgWpLPgWp/QBv5xLuXx0Hgn8FPs2DYvV+0zwAj1/9UlTzoNeYuZdcWQKk0
Uo4z2lxe0Ckm+36ZJNTWNdKc49BV5tKtSdxAZZ/BAAGK7IBoJly49gGB22lRQ222h/NINCmujGCS
ngXzwSAWO6qwTH5HP/u/Ntods3HSlU7RSh9gHxIYoZOOwklOUAj2D6P4Uw1cG5V/EbhE4qbenay3
etHCWYbEmFBS5I9P1HZnYQgAhfOCztoJ0+FU6VtnonsYGhNORQ3DNnecC0TTnFmpXiyUjrcc/H35
Z2Kz5xfNbBHcsWOPS4KYyPrnNgseR0HKSCfM5K2k+w4YgmTjmmPmEBD8RFom65BDRCjGbdblQcVN
eA0cnk+1DoT53ydp2rYhpGH/60nyu/DBHhQbU86dB8hbAq+CbXqCocq3DAS/Fk9837MywFHW64Wn
ExBbQHw38U/BHwuiIXNW9bWJwf03jyS8RkKN6utnx9xdr13sbtQAysJ/sF8Is4N8KfAnrlI2vSPA
OLUc9E7Vp4wB1gHWD6W/7bXAET4ENw3JEyrm1cVRFCLVq2skAmLN/Jxm32AAg4E8Ks1mfSY7fF0r
+C+AMhDhexe+oD9yS00ID+qqIRSpWyT2xjxrchJ3BRxAcv/fPCO0pYqcnKfCerIhhqyuKGbYJm7x
g+gbr9ccPJhAmVzWf5KXfLOJttz5qc1/im5i7fPlbS1M8bfSziC3hWD3CTw7uerGzP8LTDhjounO
6FZX/dhqXhBODRS2nk5H6CaEx86Rae7Q3qfBfMIXNzkIfCUR26HP4P8H+C5Uj9/2aztj4YvtzxtE
2r8NrrcTMpdXuSu3LfZ50kLZcEENFudcuxY2T6ajJmACISIOQD8cra85aovKRJ/+BGC21N9avY/h
VHOhO831aQdX/mHY3tDCp9wWE815ojdK26MajdHs+PlLDZ78wV1ZBEHnBsWLQfueaWg5MXR9bxMz
EKrISNK87fRG0SPtD1gu4S9uMd3iGx5+240X0z7o6Qw0+Wfe7WT5I5rny1z2hZGKi+zjrpHZgDPc
n+g0Fp/Dkz1lfjUGfH7sDIzeL7itYhWi1lIwhSJQR0omDK9DNrxCsL/wCmPU8mURN92tM5KDN3hw
F6Z1+/xtzLgwqkD50FDDyXLi+3JBMCAl62jvEaQvo/SbdtzhgYv5gRLfw0OC9XTEHK1vWBDsiLS5
yaEO4Zd904D8METUVJ0vZ3n/hONpDkkwKz9aRDn1BGeunyJr1p3dKxxQmHZaQaRUeHD+Ggsatnll
PnqSRJKEk8mGuPTNxFxJIqPMwGguASnD3sJWzck0JAis2BrL+EY2YCYvOn7BopyWlnLNST8hn4qx
oYbRYWkml/gslWgRS8727nf8vqpLmQSvf9DKVmg9tj6D+Ptt47O4zJQmceY2wuZKLUfpv3wlMVKB
AMTCZFR+YsF4VKfp155CsQDSJmiStQ/xFgg1RNKBJ2hLbR5+65quOd/9odK49GOUNMj4VC+S60wx
2ir4knq3uktOfgFm25yBPBBsgr0oiPwPJ9NlIaOSrWLpqDQG+pXciqrbYYl7KUbEAQa7ZO+nzKSC
GRGuq9cooPrjfRlNed9DOF7QybChS+iIkIj5jju3zOcVeiaUlVX4QPUlAJ753fp5n9dz0ULLOkui
Mj3hjTT7/uYhE68kfkhIf3KHmlZCJAOhSYyEgKFRohJ97+CBkWBxABG0b1iRC9MnMh7cQ+uNPDxN
ZFJ6m7LDz0Y+KgQYCuAYaPpMnI9uYV/WanuLrdmBN79UsJSeKOseW83WE9sxukZ/i0VYgoF4DOvL
gxkYXNt3ue+60bCSqQocQzuy7BPEz3KB+2ACo2qLMuTZ+bhQkCjeEuOXXo/EjLNAFk8DfT1r6Dfv
S02vFup6/S8lkJhkKcl1pD5PNIxlFQ09qdrWVJtvrFfnn/fwgyJYblsmPbFBcbvehTJWM7Io00nW
SAFnkuhbK1DOcE879/nRb7VMSz2MIp2kuy7a02JVc1Ax8Ixhm/Bx1ttU9LluDzwlnR+z0q7gimPC
0QTJaS3KqYpC0CjKohBdtlcMYvHjUvYcJW6EUSTHsp61ZlvKwGf3PgltDfJOfHSR7cBpJVSwDbaL
vlVgtdpv4cnCDAeMrG9lJYWmwBoUkE5wSQXQut/8RAxkyn+ywq5EgIvlvb2MbOrvAGr4jFZAIvG2
7tpzG8ZGCPL2/9TF7HX8xS1GwLJSU5+D3fV5OxkaEB+wooDdFMZ7cQHF2FG2m68czqBtW4+unBQP
HUju8CnfZLpp8ykxcm+UaDpdhKmm/IboZe8cjb6kOeTC/yqOhqvPED6vGfxkxIEhvicpA42hmkPB
VxQtcdVv2MXvPLdEKtCy9HVmoa7CU5NyMq8JumNPDsNG95JDRTnhmWHp+EDaauCe7l9Cla30mMdE
HUQroKeSZFJMsIiHAk97TyfHvD34m0fDu9BbLxF6wyE5XQ1ONSXxXQFf9S/9NzaRIHzJ9QMkPreB
q79IfyLWANubC8xYQ62OSK2OxcKfdz90DaLrG5dUQ7B7IlKz0TbKrs+3yaVENukQlbjOWh9bR448
NhfQOjMfsEROZktdxtu7I5aN6iWuniPa6FsdFSsz2LAkbeKx+DdbTUnZHsvSlO3L9U0QEoYgr+Bd
5PxdFGmtTY9dPUL7CTwam88pyURwRs6evgWOU4FunbKERgnRElbzR77EspfJWvIoLuHi4VIe/YBt
FryIleT8VV+dINwev4tux1qdZq3pctxfgWqO8mvTDhcX5ZwC6BLglb7TvR4FGSgtoILjGMHY9f0x
rNeycMmm7XMwrRXAkjjhuhRxBgfg4WDRK6LumzHTIyviuhWF2EDP8T/KXIiBSPC3m8XpDiHEJQLs
Nb0PVhQGVBRFX7vegQLTAgTrD0wFgoW4qdnEwOceeFo0mznpiIPmXsrqPyky32ACLuNZURKc1N+/
ifwJZgLiA7GQDxHyaNVpZ6yLbaLbB53Ejyx7Wbs1wRl5UlkNgoyK5ImXETdh9OldAVmnfUpn1+jf
Yi279XHP1iIhCQdFHPb+3XSMuHC+1ZcBDoPdVKHvZZynsfb4cbOjIZU45MfLc4qJ3c5NQ9Cu4rKt
1tLK6HNtRsjs3gzjJvmE3qTj4UiOPo6SL+3HRGIsGxCn7tTEeYPHOvbqFLt1TbZQIRfUKoZvtQ81
aQv79MhlASlu9NRseyjOaEhcNtYyXnrVI6PqNX21dxGlwF2DDhEIWRlBUQynTzJisG4z/S5uWtwY
dpJWAZSvyqD7Nf4Dout8QeXKGstwDBMMeeCcwejp94ul1/lAQLAXYELm2G4vq4ntoz4bXCiIlbj0
4KF5LXhNfPKHk+URMhCEDd+K5Bk9Ck2bpcvjJT6iyh2bf6WSRzLEjF5SAZkubfNXFg4cmfanKa2l
eEVHqD5EL57kR1YiLlzA5jxMcSsySoJ0YLOMsUNn10vCOCRdpGdiWH2YTrhp5lHCdI20CQaipyvX
IkREDIjvldBxMZa3PhNS0FksTURCxiGQ5FLN2qRt4Yy7tZhNnBwb1z/G1KfS2bED9acicPvCdwPx
huh53fH0034lrs2gMR3neYE0ctyCIpD8quRkwnWgq99qrmg25gfAnPAlNGvqqQLw9fGruR3aXHfm
bYz3vtUkCXWKBOJ/VL67eU9lVKnhamaEOzWel/vYie1o7eF53/ykJMzbMKYm5cRpapxGJb8KmW2M
4GlKm7PK6UwlLlcY12aHnqr2JDJUZdyoUWShTHJXdT1z1GVdsjClk90pYKZIIto+7T5V/cQB4GIg
PxgExM+XKFtuX70BZNAcZf6l+D+VXenQQaPwcanF1zUvBn+k+yF7bL2fekdZd120zUNZADqGiuWP
wudwzIgtRbOOzBXT8dVoPG1UTc0b89mjxQKICmPZ5D9Au+ym41yHVFxVmymeE3YTb7WgZ1XCNMla
Ro5gaTrnNCroI+IpXldsNdUTJY5ERYmikclHEjVBK1FFHVe3IaG2hbFXly3G7gScxOtdd8jhRLXH
OB2b8shQS6EhSYcTUMCqNDVyFUwIPPvL22hifEw8FsSw7O/NOw2Daaf60vfR8uGpD4BkdsIz2Q5l
Z3UAgkTDDFfu8tE18rGLrVDkS3ehUnbSfDVsk7Y/lSwSuXy91foqUfTLuyHLGuly1d07bDBPAYkI
7p3cNWiXIK2aPPIVhQPU28E3zBbqs1U6yeZbpp2dymuf0ar6wl/U3jCMJ80Ywe5W+q+Lh8bzkAnf
uJ+uRu4Cg5hirnTSaZPqyVKJ+c1Ag4P4JODgcPyiY62G8SisToYWbiiY/Gc0sTNqVMvXj3ZrsdF7
j8gwUIfHK0A1xRA948KYk2eO69uk3yke7zDRXSOEOQ2xWF3pud0wnEyxXtSshkR89uiQV+QiVrYA
QvR4eFwlHtoOYfK++9hLJqfoYrJbpFEfgH0pp5jegy33Invec9QbIZNv/ScJrTIto2fpXI05I9VO
kcDLcg15q3+/qCpvIsqNdyVspBmdBSP2i+VPsCWhi9nuvTeo7faMOdQWu12wgotEyxuw8/niD5E6
e1mV8B+yh7wxDY5QZlQYVwIIhFYrCBQ5Q9F7xtrX9/jvlFHDXdlEsGBGFj5Jl7W4BM4PM2H4ygZy
J6M6FiDUUE9xm5m02UqOx38sku2MKzdSUVNJFDuBppgchnf5/F+1uoMpmrsx1Ah+XIsjgzCTo5Ge
FdmqDNrwR6JvvDaMhryKXrKQ6UMpW/zfe0/GWlTeuWxv4b/OwzFBLMr1m2/SxaCWy5JNFucLGEY1
cSg8RksAb5CKPh/u8LEr17NwytI5pRK+0OCILlDe6uJIADchB2oTiXhVukw0cDRxwr0yNqdeuC0L
DuaT5FawHFhixt25B1R7HAscygH2+OTbHVMZTIYTLAmBJ2nYs+IRJ2Cn57zeAmHFUnOQ7Ir584uI
Kor7cC7n64KpmSAD2Qpdco1Z8MB2+OqZG8+lymFo+Dtm3+NAhBiwkhK3nH7DtS3UTC9Cxt9rO7JK
SpSkX48cE3eHu9aEzLpc21lVkTX35LEmWAlaIhOx0ftw3OAGb5iY7JzY3j2sioG+v/XwVWEqi33y
LiEp3cgRbmoMKVXJs8ZYMwpLgNXMig1iu1b/nyIk9NUvvj6TRFdd6A+3TBuynMBPiKF4lu8zrajJ
sW7YeqDtRheFe22m3c8EI8djQk28lCo64oOrbqeebWRQ6IiYvufmKOwNBejvhgGc8W85UfNARnE2
nKEWYRoBKQxyoO4sAba+3l8Ss5vcfiSoc/0dYOeCbS9SKimZvRqTLw0i5j2pB8+DwygLCegk1Ltc
WycJjEuVA2PmOaCPrHu1ZGOI+1/Ucbd9wbzaODm0ZqKxiT3ASwxWEPgvuTjVSUGTqgxvCDvGvqK7
0dpNl6vHhJ/E3AeUCHK+E0+/YaLqPKDlWshbWvChmwYvvOPSrtjZmiIf7lZKpz+H3nS7GxpKlbjs
f3bPBMe2vsuU4J/96+v+doFn/jFR2g/XZ6WW6Va0c/V+MgrLt2J/9rmdj+bc4Cc/Oud5wu9JXaym
SZImAIJK6NGgoN/ZoNgLuMi5JlUCgcc8miocM3MfWOHABX2Vd9elIyiR3eTJtiLSJKEfIkW6ub6I
YNJsDtIbz9VUs3XJgDjIjdePVILpN1zKGjYO0SlTIa0T4/LcCR9O3V2nUa4PbVCSia/zvsYXC36l
nZGOypk6b2ynJV4O4L3RsQVHNprjCHhDnFH1vuyP/czyEHn8Y9gsZhSkD74d4jRWjli0ifK0LW+8
9dtBSBh2l43WKXa2bea/+0npo0K/HGzISAAsnT2GrklvZ9yv6SMdZHOden9l7/1DorKdxIDsQP7a
FbAsTPCbFiOvcKtNCSTbFpf6yaYjKaLKjkRqJpTPnPLvpm/A17yIZkhKbkW9ZFWqvDP0vkCzg4cQ
nc67uqAwVSgzaANkC9U9TTJaVKrHm53+h5rWVo5E0GfuGiPVRi7vRspGPR5rh51UECb0QhDc3too
PPZptdwxmYHw/S7Cd7gdGgxL3GeZRe7LNjDpj8ActA4AaWFycMdla6KM4NAd07TtbgUcd+2mfI0s
FkGQW4KXBURB7Usbq5zqkVN+cz9OJyhCCM5PHhNXHNB11WoI7ruoMgnnDcgenIeoObLAU7RhU640
d97/IBCoc/Gkq+vUtKOBM6ci3TG4uQUvd+dQElGyWClgVtuJPTUGToCplWxsZnDveK4ERRAeCW9e
Vt30IVRVNj7zPsGOG6hLPwCGOgoJuZpoLBrvIWWpbBRF8cp0V1NXUjdI9ZJrDJ07a+SdsiGvjqRf
n/8Zf4g1BvXEUuYHpLpL49yb4LqcXjgYUGP9OjQZmE2vtAqqgKRyYEs3iSG1CEbo7tM49BTRMiqV
NorU71BImacBj3mIEeJHFAfqpT+xhWn+YBS+9bordNZzlHAt36R6nSAUyWL8K001ZccXlC9WWRi0
8qvr0GDbOthvovJ11cXgX/RscmxjPKNvBpYNbFWqu3gd6jBGdpiXRO87+Y+dQim+kbqhCeTd4IXT
U++XwNFkONHlsBJspIxMC3fmjoHWXtvpmdE56WwFVufTJXEQ6Sv/DACgGEk2h0Kfp//MNZKP8d0R
8NgyIkgZK8l/kSlzREIs42dQwjoMX+MfOgs7NCOaJMSfs9L4ro1QQcGToY9P+l80ZmVjjkV1YJu4
JyGNsgxWeovjIxHdXgM1iEukpoUb82ur2a288x2NYhm7jNQFHlHxaTEgFLWCNUdaKmApklA2m803
9onULNJX6IozePE+fmnZ2l/axSlWvIPtiaw50S5uHggGd7I84z3Ns1r7zEpQpQhiavgwbhme68sE
JjY/7ncGQf69Hu8rF6+HAF4S1PsjcDNvs6Hpia0v76lZEr1rbH7yUGuNCpjc3kYjo0joDmLTY5be
nipM/GTAPRsNpqx6fQ+0v/aijqIO0rOSNqaf+JcHQ/RAzCqNmTNuEd4DNG5Ez2zngYRet7rDDS81
70kVG/DCodiCT4/iM8u+ucecWFnWwLVQ0h2ck2Ld4p5WJSaWvGB+H+HO0xrHSA/L/idGXc+20Fjs
ZC3qDEzkwMEhOXRiOl8xWGclyOcGmgj9+9C0DTh1/tXoT7+2eM/tx2nqY9ZvaSV8ov/lFjNnBzbG
GH23/eXhcvotL8V7pXc1QDPr0exE9yO1DkVRazfhy/BlKRaZ2Qj3ygf2OYIUs5G6vJXAIVec4/Cx
MCK28ATTqslBfsYNd18zOywx7D3n8t2HsbPK/3PA8uPknOMAi1EtKEi+puOknhZ3LowH3j8YkV0G
4h/ETsxASMXCGkAQa/wS5BG7gfRMT7t3kYsxBwT5gCxXuVTZ3IiJWQmagD/M12fDegA2hwYKjVra
UGKqhH/CR4f7iiKpRUemXEn38mZxklEv6loZi+S8OeqNFSvJdMpaU8DgH4q5tHKaoDDusns70xik
nWz+b7S53ngszaYpGis5kf6vtVMz+6LIK1WAalC1Rgmn7L/sYI1GAewKKN/7S0RZPyOsaZ+wrNUs
uNJEuXet/JzJJBnUra5H8NacnBcHv6wGe3zwuvBvY0IlXcTvaahZh+uNSNZu+0SwD/NL9h2ztuqV
+JIIrBpw11teF+RySKZ+3Yg1ruRiPSp/LzdZh2jlLFz0U36iGTFiCkPMmN5WcUvh6otqeX0eVgZH
JlefRYTdNX+OAf70JiNaLsxgrwdNlqUsSk/bgySVsMJtNpeG0CpUOuJHmaYDo6bJrZVjigfseqir
nwxPqmiBW/q5RqQJLuNT427aF6kylCboWy58Vohfvu8U5DpwVoFuEPk4anvI4IxfEUU6N0azmjjY
KsWH7X7gk+SwnYD99k7TvxGz/FvjaT4gaVGAcDlafu9AiXJX4OgmUyPM4JuYIL27cJaSfDLOUj34
1t7onyeHcO3Ro+MO8AWDphaM/g+PiFVxSZwZMSWx/gdRJN4MRSMOhWyhEKeWgkr2Q/obctU26CPE
+WqKCnWs6PU/vwR0B3SsI7t9skHiCQDspnSzecUeSsdaKEQR9Egj0/P+6QiWdBx+KXxiZpO7efP7
VY1U0/dHrqLCgTH2vR9Xz/SbitMrMJX0LVMsDf+OYFiTePam6KAktsjxworVuFGtZdvhjqdkYQGr
tbNEU+4n2ZC9nfCLKnAVoso+aavdxjdS37MTVahBPTKNWT5zdEIrdsDUl9uyixPJihuArRzGYQIa
SSdUrpX4AdXnF7pMAcCscb1C7EOIMO9cyA+vaqUP+Yb2eKmP856eYkaXqRPYzJwpE4oZGdxNHX9t
yE3pQ7Hwu5MO7qS47AWgRYU1UVjCd0Z3ZdbW78sxuTD/chzKZOmYd0G2rgnOAswsIttwoPfrJ6XB
NsAtdlwws4atdSOk+bQUSWUtA4T9xeZPG3CqWSKIESZ6nSdHT25hrz2Z3rrBIqObaSJbU3+QVJUX
g8fM5QaTQwVAvgI8jRltPc37GX2L/sS2XCkGUYeYbdjSN4SzkevqLKwwgSLFa5/RdT1IDTqQGfHe
/9gr4anV6+DdwHDQMVc2XNMkgfsR2oMCJ/uW+UYd1tvrWsNlq2MtIEq2VdMp8ktK0liC1MJ/OP5K
2mR8B4Cf7E3JtNTZLr6lsmiJWMZvH0F2m4J89BmKk+Oaf60VAcvHUgV6o7nGYAWt9lpSOTCMWtHL
Yw5qfkIPGN8ddeJ4YYOpg31wVgpXTl9kdfKaBZQozsuhaupLYpnHjq6jQ3XqCXmw6Q37iuxSXLks
Vuzdq1HWTwUz4fDbgSGLYkn6qavO/pLBOIB4iZdYh1ZXO5P82HjkgUAu8RRW86qsasjNSDp72jxo
n161/fquGq8cfmiO1QDGlJMrFP0rnPTMcRJZhbnu8DR37zVlRBZOJobNPeMh5BSoQ1HRTZqY0Hf8
+k98S5oqKefIuWtbastPp7W1aYXii+rHPPE/VglaEAYDEbPGPpLpssb/xegf7rtQQAYYH36iakmR
HkZrPObAmtZATHkJKp10iY4MZOZhwUcP2SBRHb/RE4rfBb9PEGKctUnulc8L+d1X/zI5YSniqSDQ
6bAsIgwcArzK77TUA11wCOm97QTw93s9mYQ0IsMMS9yHjNVMrJ58vevpOvQuceCjqKO+tc/hG7xQ
E0T2qeHijyQoEGLYS7KEhCnpAHzctRRIstcjSklcfdtUdmhGi9NEC8+VINorLmAzcIDHMwsFGoku
AtWTZYf7rrBi9XvqNHKx88ABwfDzKK7+VuFnKxMwbWCzF1xEu3c4WAmVa+2qv9JnAVd4k85j/cjV
pocsdGzjfdhS/08lXzsoxwzRIsk5SlG8A7M4uhLE8QOrXAmNEQSiHEWJARd616cd5rNx/3vtw3zp
Nbi6uygAwPjTxNlrPUsGQfXHoJmcjSy0UEsOzGBtbbx+ikCwjs4mHO8cW8Sq9mzQ2/Tek7lmmuGl
FtuGbMvg236lhTWa0kC5LHIyR5reEQa9+s7wfK3hMrApSeU+mquEc/J5/0g36wU+rxTo249ovTGT
7MJuvD/v1jKKIVKV5JQDPFjoQ/BOdBF3aSsEWEujPduZbz3ceXZ3BUb9V2dOkwhBPri8iDe6cuXF
MNFXpM/80jvnQ+7g8e+SRZHf2a6cWgDL7oUxKqYEQoQjJ4Z8GDxQFr8E7UKHP32TVGdpvn4I8Ea+
/9Hv4DdlBLftYe8Buwm0fTzAjEWykF3sIJChTgrntEmGvCmA9i4+suvHeIPu35oDWm3+WgnzUp0R
JuNDhrYIWLDENfZDcUszDfELp4EQEHmvaYi1WD5pDzzcd1Cw6Wagl9Tkx9QhiA+FMQB34HdZBsKT
eVEQeWZfk5f+gYR+JwxsQxmsp6FGG6t71HHzgAWBJcIQyapUJ57OGfW5FsKAMDsrFrd0S89FQk3+
D64/LCuZeh6Hccf7OWXN40nQVk9zgiKEbmiwghnriL/JOtMiLvlby772l7GBgawjX0meepNg4/Gv
OsbsO98qau63tLUP5A2gZhjJHaG6X14+tDS91TWSYH76UuGHEobIg4EUKyEl1XGfELuxQkmge9H1
NOv53CcEAjFhvCLrUzIiiCdwONlMItdZ8FNZq489uCJeSXSUezFyRjD0PrqFFz9+q10G18VMyNt6
tFmYldZhJQ+CtI2fPSDM7ugwzIRobwYO6HjhTjRTndtR79K9eGvu6EHKNvwJFk9sT6jQqYr3bWK9
qT4lt4yAnuUeVmFIJuVD6SAdIN8AuKfee2GwrPHcB67HcQXsYlogRVPrHwYRYFVG+hfyphaMIVJc
CJf1QKGOjBsfFu6xVelrc7jbUyEG1GJui0Vk63Y0E+8PXQ+1FOpFkeJbginmlm7xqZuScQjPHYba
asYd7vEDqqhZGahjrQ8yf00k/11d/BaJboRuR+I9hu8exz7zeHA+HfKkVA1r7PIBPxUmLOHEFB4Q
twp0QPnIYbA8mBCsRps3kLWkQpOWGJGJ5xZ5kO82g2LqI8m+bUbuS1aTOzNuLgXh5V0S/ISPxYNf
bIvAPPvA+ebYbN/3LaSSlp77paSleMvp3/LOHpRcYKCLuumEaf9/QGTd2tmzptQiQA4wI/pGKWVS
yyBw0gPs0QLAIqKv/IT71NvTN9hcejBWrON2In3DIsEpeVhasybsPkr2POtNlR0SrZmtU7OSV50r
4N8lLnjQ++8wehv1CFyBZRkRx7eXbrgHNDL4McYZvtSkO/8wAU9za19ip7Pzbw/RVFqrWLxyDs8r
Uwe3NsS11KsV+Gvklne7ZmX5G9AbZwsjwGDvzORxwtnkOBkCqFUWc4LdqXyzAhs3r+mJtIVh8cn2
NlTBMCS7CfLODentU2+TEOiz1M7Bc49TzZm3uWDTsp7otQAk+uWH7GqErTNARxzFB/OImzDGWud8
QQJZRkDvbtSBZdj/72iwFhEMuG5kktwzG5rzF75NhFWJP/2bbzuER+HgLxh4rbYMuJ2FdNfoFPyp
CjVJxIxPK8lRVhCvk4qyDV5rXvKMNsstrX/45OFLrfRKCqHsmZ62AIEC9kruS8JO9zBQ4M9rfmvY
uT81N93sOaiuF9Ow1/qEie7MmwDKKtaxDn9y3FpfkdL6uMUYZNCC8Cw/SyFDjjBQClA3BlE2qcOp
ai/fSZuGdq6Ge0NE72deKXlbqJteikDn9iPkGDIbzIlIYgCGf5dF+8LrrwnZqGkMofFx7+CfmlwO
LrwLXWHaP7qF/dnCdykaAcg0b8UssuZGIqU8k/BVpYREbA8vqZvO5keRxcVvqMn19mieEMJbHYma
UtiyiV2s26F0K83Omj5QbrwGPyNxy19Za9bm62WaoyJOlVhPxA5t/IG7FCjDBCdWDFqolDSgZCfL
byP/5oScBYhsoYUo9XhLu4tgN3Aa+ToMkMXV42qEbKIal7tSqs0W8O8HmGfaangYH/Ke4ExkXDBk
NWvLwq/i3VSKPtEWwkShDyjVXAJM+DmKLxRFachW2MBwe3d1X9K/DGk+9lqmn5058hLoJnAq1pZ4
2cEjGNA1Acoki11kEUvEg25coe9/hfghyzYazDtLdXWJcIjveL5oUYHon9Hp7YlECzrYUYBgGqiV
rFZ0MD2LHDHv1NKIIvDyC5QbPNotUqwpCzBw/KcnUefTvdeyLv+XAPFaEiCsbqhnHeIjY207u4hn
kGMfWSqTFdajxb9QSnnVqSTSywnAo/qcdBKcsnfD5jCJovW/oQjBsN5g6H0/3dAFuqahWJrzJKyK
qrk2Cf15VfHIvzwxnGmNiSVeldTAjZUfam98FbE95ICj99IHdGDNJFG0EqPkix/fWNkE5N8OPgvQ
wTunYROp9vfMVFl3KUW0eIAx4RhcDDbYfKK3M0Jnse8ibCO90rvPmiUZCGyPbcamxfFOAEUJIX/I
u5LyrWjUQCfnxPTyllfL5/hg59tUUlsdyxq8qpxNXtTbHzI24u0I/TPmISV6YNr+YgJZXe71tDzv
6OlrIQmWhfvQhjAN1IMXG4PYxXlv7u0RsdbXxyo+jC/BvUDCRRA0WM1ZcqkGOuRA0/lY5OwABNw4
Jeu28uvnPWWrq2kdq8LzwgTr/zeg7emZgiubwjUtKC6rCIvxhFCxlZU5vn78dlYxeLxHxlnIRrN3
2fYmMlVgQyvJR66xQN24A3EcuYqhcJoynTQNiycnE35mkgLM+RCKPVQ8WyNevAzONmRgAFFCg4LZ
+14ZLk2weYQ7qdEIffSr/0dbww96+56mCd1JFujPlVzCGbY1V78eaoh4YKw6VZaZxLe34PlBgJQd
gSCOGYLJWcfs1vlIbiQBZ/c/anOgeILfQ+UKw/yII6NGGUvDjocR3SYePB1Gv0uQ1LIOBB8AUnX3
oWXzt6F4geEC47LIP3uq5xfqMdVGMr9GG5wsPPb9KQlXYLoGtz1DwiYwjK5hXDX73ojGDBYBezOe
1MAMCNlzscy/mpN9adQaCgPr87XkLh4scjPIZoiBSIdG+PkUXnpRUaLGNgMnbg8I4GvS0i8exg5l
DyL9y4Xyu8pI+0p1ZpljOMKCtP8cUokBUL6zqmCQkDukWXSTQFQaY0Lsngvrf7hbfLikoq56mb69
UK5LtH5V71+p4ZaZRIv173vzJ8Rcgt7cTlROB8HS4VL+A5xPQUpfZez/VC1Kr+4A006zxI99VqFa
s4DBy1z8I9H7iAEhifbeekSCxaYkwz2XS4/GH+xd+00BkO+gNsKzWTYYkpuuCrvOk9my5paMMs8U
L2WQ/dQZZ/n+SaRs5FkwH0ZvO6YyfJamkOlNAdZG+SbpOtT44jxwD9UoyFPKqkDgnTY0Imc64rwd
0P4l1t6bRLqC6DAbC0lW90Blo3HZwSIXMzFQ8xA3QxX8udcwJjPNaK3DVF5jfkXleQb8HiRKcMlb
TLniFUlCg84OwhQPFG05PJNhp27wU1TUmD5RjRZmpoQGbC4zAqjbxjicx1cY7ZyE+/mozvmVA8sc
8f4nCqgHWerWha8PeDoCR7hWojeERmAi6zcP/ldthxGQzGNmRDCjwIr0Vo9JV3u9hFDFcmD7Q8oz
imkk/BwsAwPRyOZYcW3W2dXDFDuICcYqQIOaq8ucAZ7aHMG1MxKTX7t3L9yTCnQC/eLY3p414Zd/
0GYaxToTVe98Q3aEYT6qUbkGpd2PYi8jswysBTibizVfETYUtrz0RLj4urQoKgxDExrx8y1jvuKe
thbBegVzbBebslYcEzA8g+XIBpO2QY13B1hlMoaAGmvSryt60H99bU+l0CFuSXGuSYzNVgOPmlQr
LSF4DppzuUzRmdLoNUwSqkFhMfL2Epec+9BH8D4qFhyImhV7FW7q7gvity0m9BADUNqZhNh6jYAe
ueAvD859UwwtQEO5jR4iCfJ+QcQa8ChcxbYlthnpCPxUclVKtLZelDf+QSY4hqMboPVa/CIs3kfT
44CuqAwz0EZaXML80xCWDuQrlCMbKVFDTZY4WKVQ1hojI4ZEyc9c5u1metpMdquqKu/ntmrtLGcn
mG2CrknlvfsB8k2Ycr3s/LhBVYLcZlUQ/nLjtpsanNw5fXosulAM39zwwlNiVyAoamFqSKrG4hW6
YSjoKczXPrWg6tkEUCBk2L1Mslq/gxOMXE/li+4o5ySRyLnbMgefeFDYfWqvOZkFZn3712JJ//Ni
EF/LMK7zTfyth+xi9+15kt8jtmiyXv/G++xpZ6iEkqicjygGQ6D93b1dRnxu+4IcN3hE4F3ZxWry
13zN57OweXLK46bcuQS877hQh1oo6/+c067g5cXTJ/Rt8vP5A1QZtl39rVC7vDFH6OI4W8th1Z+y
dfWMR15FFvcdZLY1D6iUeHzSC+57LiyhzTeo30J6W1mvL9nQmETCMD+q8QgejXN3rxvv1FirN1aH
uPRYGYPe/d7HLTkTgDxrfL5zjK9b0BTAtFgUSMtEssFcnEiX94Yc3RwL11H1P0Y+kccUmp2ADVjV
B0+YvJ0xkSzkjX8Z0nw4kBcDpO33lHJLpDfBzzNOUGtFE948LC3OoQIUtMtr7S5lp17t7yHg0jR0
JTnR2XWgxNZj+wRep/T8bxG8AUnZyHz8Z5lnN9LOJF3r/5m4YQHcGNNufGD4IUFdFgK788kLCDmq
OCQDjXD/8XGUdC4ZGoek14uqnMkDFgZjXSFBxjlBDxaG0GAXp+MnC1zvzEbSPbycMv+lJhojd0rr
UVdSofFFMGI3K4vBRbkyahXBqC3rIJmm7mQIFXqd19lHPEoktPZZGwd8rczKDFSeMKcZ0tNJ1iDr
c13orOB/7XzS7mqdDNfy5M9D+01eYZNgGCNolClywGtOX0aWi94nqWFb7BUIzqC4oE/gApyF7CZ0
xAEd3+rr+fJxNQJcLbdHf/A/iBfON/zbH/RmXzOU548blfB+GDviSxfwAqz11r0g0HCNBBDvwav5
hi1Pg2s5mwftsj0ck2vASTCnJbbBE2ndHYwtrwbZp8EbECDKqOlNqm+h5SCqVILQRLcZA+GJtgtL
zN8I39rTo6hlE++Z1Y+TUA0fZlHWcD5wjSCPbQoc/wpTxwLy2vM/nSFJOK5Mx03eAJh+zxkrH4FS
Y8bi8Xh4HqDWUXSL+IVLjqAtWaj9KlsImmcY2XfUVhTcFWmiDg/XtJ2/6iZRyEOc1e4munj88RM0
kFW8yWC/gP/pllcLZndDjbdgq5wcsDbc3A8T3wKIBRd80Q2MEhx1kl/3vxu0ghl+0NBXa7UVWzPz
EDeTO7GfvWh70JC2BWzWA3s55L7gtys9xTPU5EfGLij901hu7ssYJRqMp/xVFKAuar5/22oVYAEI
EUoxiJOwGwXHm+cfCotVDuSnnEXfnbf1zbcgUBvFEhANVJIMp2rEI26kjkI54rYvtBmZsvgCe82c
8k3cZsxZ1kp1Q3mBBDK+TpSvaxlL03m2T1BlWWgHyaFw+O1hwnqhvOoclu824H84Dmkq8TBOStHk
JSlR8iAH4f+vFh6KRku2UifvWlKkIcBaCsr9sjYZXr0nMWCnMQiAEkBkPj8OeDH2WjXaVMOXGR0v
/R8DD0F+Dvovh09YJmqGOOSu1gRBwvW5g8KTyi/R8w07Sr1kTAFf5+AJr2ZK5udGasXcZTOgAcw0
roqglklwuJmRCLGiqRSbFLiwhScmjjJb/JU0IcShfIQ0J67fBVy2lXOWTaKKcersdY8X2caUh3iD
6SbOLXSDeNqXSIRCedzKCpArXMpGKTzHlCM9Ghl1D9QTtrGUah0NVZlXftga2eSAiS0FUU2jJ+oi
WsunqRVlp9Mb94DnunY0+brEtI5aDUEaX2i5ecgl8i8YHxHMp9hMSLa5pDwaa1tquAk+J1VpxRyh
bKut9RGbpkq2YJpwBbr9TX81oB2OO8JgQTTpc/VQVYNvGbSyTQiGrbe1G5DkEbixcsbzeY5Otnfj
zwXAGNk61WfqExkykQPYwk2H/aiIN9uGy/CfuBLtYJeD+MyfatZtEjF1PKkwPww2WEYXBpiI9Q6N
TpzJBh+LNANw5ZMWF2+4ToREyJzsW8g5RGAn5OTjilR5bAD4DuK2ozNrfHOR+2UXZOIVijXG9+au
7FBN6FAQam0blMkT1rYUCv8wabopKvY/h1TtH6WfQMwDSvllYzvzbz5KBlK58/5cG3LpLI2s3zm0
zEdeZEDywJ+qQt12eTzWaU+/jOX736QDFLF4rnBUJSNurIsWxZp9BLy61xCO+oVjhRzfIB2P4Txb
jqvSHGxQaQUJa0ambDL5xmWZmgAK+hAmZ9vuA3OIZdWSoxjryZ5lwZ1UcKTpv9YmLNHpUHVd6gjc
Kmi2OliY9Uyvlll4OAcIR6R5b8W0XGgiu6hAfHLcr8Y1ZRhyguMyqwJIWbtmZGB3O8sEr8kSucs3
AUWHgOG/ZfWdLEe5wDR9dRQTgHJFkJW7PJoeZKDYESLnAnHYdn3vuU/o0cNQjZLPW8T2nU4qG3WG
OYWfQmuVBWOdpXURA5Vzm5Jku0xuzK8O3tovoki09WFRl+7zdafYAgErLobW58nzgGLWqC8EZAlm
XR4SkcT88dc3AWChzjITSkvGnDdpu7y67ik1dxvulIHSDjI435UzFahZlg4z9UpcmhcbtTRjMDX9
/NkbRf2AQxFCxMCw5BjEV31AzePGTyoitcQt8uI+5B5zyNBYeCU3RzNAi1CbEQEX+IqIVgWzFK/d
P/NLvIOkROEj4x5NRBZ0XTMGyouAVfX5xXm3nsawCDH7cqp//dH1QE+ls5gt6EIOnbHTfiHoELIm
A8J4BciSJPWeutoh/YnU0RkjFLlywry/O5k8UEgvp+gpEiC3yl7ewxvp9LfkLosKfbZrIgTeYLDi
8kiZsK5ovjzKBmGil+7WIk5khNevnufQN3U1lsIX4PA7BUW80UsZ6KfJR67aQAixJVpwuVz7GAlE
lPy6a6zhqFB6zFObVZspYG1IG4ZmLOiIwUOFHjwyAbv/wmJZfis9OD4omjQvfue8VR9I4hRY37Mt
Xjm5Cp1WmZ+6YT+S8biP2DbFOPX5OicrnwiE2l9X1P7cf/wv6L+PHAVGuPsLUQn8nQFq/J1ybkKl
kZpfq7H7iwXmKl2WU1qk1TvfbOYPAnpuVkaY0y+0avj+Oyh0Ic+ixqUE3qOsBrPLtRNk/WQD6sSZ
mdrhs/Ajdtv0ELpsj6qfTD+0rEIfz6409IYSy5n8i2Pzs3WdIMO/mDCP7+To2HTuvZTIN+uP3lIW
w534/Dyo6T6uBarw04wNJWgjtZAtcACTANtvzljGwZIWiJxTwGllDJda/GhznZmO1/dV8fNA3U1i
e26qiKhWd5mDTg5jrBjTsF2fHWavJgWydlh7r5oOKp3sWQXtk0enSI3DRrhYztnwU2LmJv/Xe/Jd
axtzsdAy4Alan2t4RRonOHK7S5g8mtxYAN6Z/+bLgwas1yEU/6mkFomkQNKxVcraOQQIlXYWhDSl
IiWvfZMVxr7qIfGFScB5u0wHnwmGsIrsJ6kHrVZwsa9uiwXYdNlVQwMbWEPp96uI5XpJ+w494O+s
yrn7MPnUZwccGh1Dxw9gLYXOivPvd3/igtu7hu4IU75bhp+LV+CBsj/Z/6RUYSNmOc8V96GbQW1n
6pBNXEhBcYwjBawP/q/UoXygTfFzRfLLkRQEhssSvMCxsjZeJxVfD39UqaR2ZndA0ot4MFdqxwDP
d0Zz+TuJk4HQUgGGeP6aW9O/lQCNK7RTKwR+8BufnR0QQCuzNBx0OWgAEqAzh7008hxg0BWTHwuk
j7AunUL7ADse+2V4fqwfgh1Pt0kZaehBt03kp97MwPbfRfvI9+pZJkhRft9O5zxPxsvL592tQdeZ
q8urUkbttBV9D27+GQ3rnu2/sMxUaCfe4ANTvnbvCJ/l0oZagdeUHNvZQ0IUziQ4KgQSdGhjlhPp
9DJHtYdenMd3VhryHvSM8LC35G5CTTWYW/t3s8USbYr49PEUSUxJFlqfT4RYkRWh7UecnzVR1BiY
yKk27LtU3ZlVSRF/mMVvw+ij/7K2/4jqACo5r7L4b8kZzhYHXiyXt+RsT8gbZTi4AH/eyXOHB0Te
gb7CxZvD0Xk+duHY1E8dhIKhTPuuGqQvkh3C4yopJ4DYNHNXgBvWVipR7dWtZEpJiiaLXAw/KvqM
1aOTbGl5HWuOCBMtdDONo6Ve635GvdyMlCyfgI7YCGt2aVSIE2pbkrFGV8GlwV0PVJyuCKcTkXWN
1iARMWHO/QnlA923geLgjp+a5FTTeIYQQg/UXVwJGYAa6vd2EFo7Z7zOEghc61JKDYuU7qMsgwD+
Zv1LFFWEWbHlsBSQoPxzUS6ssKZLmaB8Sul6FrwzQ8GoptMJZ2Hy8LpqIf4gfjT5c0dPGh83CMKN
gnkSZTBNos4rulAtDb1/e8A911FEP3p1MWf8LwiX+gdmloZBmMuzfcgvcLGF3rTKq5JSRKuMTRIj
sCk/1NdkJDUv/94ExddQIOsMjdC41u3Lxn+/xcJs2i3It8tz1jrZQRlSTALaNnICU+oFtyXtqPt5
pfsTb334ipKsvU38VuqiyurAHuN4BSA26T+VY6kaR7Ib94PaauKonHOF0WbgvDVwRiJ5J1bl6WEC
svl1bx98K2+BrcxcZjLdn0L4Iro6l7DcGkBcEjl7gxsqNJ+tYYSzfCwmfvrPScaVXb3nbeoBYZTg
XXBYpZ/WXSQf1vHg2A9XVYpKbVs+yvf3ULPogcqDNFeSpS4sLvpiT3cjxdeROocLn4o+D37uTEOn
el0D88ldFY7/PODVwkKy8m1J1eMnOCzt0g+k1d+u9QHzaaUxCQzvECGBTiwZEu4Uz323vZFlw8Fq
BLv4Il7fH9FqZ786T1FqH42MJIEMJcnrG/MilhvUdhWAtpXmuPOxMlinpmSmvUgquWd/WBU2yw64
CQ8oiICkR3ywKpcTBLryquvQnzzhelY/cSPe7HUTLxKu0k/ueMpjghl1NuHXWmfAR58BM7O/6lGt
CzUHTXnNrZpLiCdaoBJ7nJP75xG2S1tsJKMpUAifIOg5LLw01kdEaWEKrFN7iAlyNn7282P8aeJW
ziAHePpto6UtPMWObV3RK0IHMXTTzjzmSDpxrUMe6O5nVv0mkHKL4l3+5qIJ12lP5tLbCd8sJIjy
02iWLuI6xvwHLr0QwiDPkpU8Mm6Ipp/PrdoIBl05KLerVYyx8piytNm/3InZBNYqGLZS3HRdLu7L
9BnizhDgaQavjF1KmvjIYsXR9TVGC2jtoqkICSfLEeFTYRsoPqdX7Kn5hRg3D0/Mkz0RkG5sSxfu
auZxkCqyyQxN1mjtTI+YrdIZA5iif22/+J+rg4dCbyHsp5XtIjCWxiKKuspCXUgufMcRAl8c0+rV
W7rPRw2R9T6Z08dr+1T+zpLH6oAEzGveTPxgjeRI56LgLz/s20amFc3v4bXvXqz8u6xYcUE7S3LJ
KAo0j7f8VHGk6JcSELDd8VV8ePV8HSEzhqWVXlAjyQjtNA0hyI5D6nPSArCrgFWT1qBslD6aK/SH
vI3W1JiC9T8D+9tq6Z0Hqd90kii2sbI/JBHHD05Pldij+54tNTWpjFZ7et3ibF5ond9xN9jLEPFT
cocKlrAMxtFUNlKXtyqoSalu3o2XnpocaCb9e+LEON5P8rDHdP8/A85XgXWxYJ/fJGEDIDABSw0t
FPJ9NiaiI2UJyB66PrGXdFckghVD0HwUS4skjWP2wL4FeSKEHkUJhBh1awgRQxHJp7Lcdy6Kpgm0
2g2GUSXZ2koBk1V1PFt0HveSMcAp4HoPeYkMGlWFV7kntqLdNqRuP360SQLTh0Caui49aHbw5HB2
6yQXUZyk8lqJvGDU9prAnMb7dk9XvqLLW8NasMpFzHpET0DEIeBUFr/6CC840Z6gwKsY71tU+/By
9w6X4KRvfXJBEwiHY2rMF4B203WaDz/+dAfJj/GaILAVdLC68AqvEINs7tU5A5s3cXt7hXueYVyk
yzGTokGiDWko0V8gTcpRyh0TebXI10Lsxzas9EPtZx9crPuEJfpm1wwa9s9+wuTppttNS3KhjO8B
IgYjYejsgSLPItG6Zs09IdCmzmqmF9NcSTSL9Q/caGGM+PrdRXssfwC6Pp+2zZi6s7r+0NAbIKSQ
D58it8U5ssmY91tdifGdOwLGgV6Xyfub+IDT8qSVsCLJsZBZKn+8STscMXH7t7bSKJ2vWTUrCOfB
OLF5svU+kBmdYiWHzgIeoNcm+v3EPJagULFqgJtK9I3ZUwggufrqMCxawiVTk5rjMO+vhvHHepEV
ewsvOOygC1024PoCJod+IsfM5umwvi6sUwkhTznAGzNNuHU1kXcJVr7a6zfS/gwbpS3hL4i8alGM
EVjKXW5cu0reehjt5tO2LtVTcSX1hpQc3vBVSJwUrimBhvk4+jO4M64JsgI9zrYteVZFicig0E7q
V1OWY+GcrHQX26h6DvQvebfsNU5uheevlK/Ve8oC+GK6jYAWTLM4ROREbvMsO4IJLc44EpS1vzrl
9qCn1SRz9A4zix7ouFTzDkeLHtcUFsweefWHfSnfITDtLJXeD6Og7hpoSMg0Y4Fy4ayZR8WPFN2E
gQArw0lgJDGxjQ4OPdRMnf6QoEfeGy9la3DfMWzwUZsFuGYwN1taFHG4w6V9tPDZzXTe8OYz28/P
9a25ofJXDsXNiHQ3brfbKQdAbZto+HWcKzA9Zex7eik+YzufwNzczp+EWHYg9jLTBM+hHSya1or2
Hjq4Hzz3/Myfp1ugqc/oOSTlsAuF1xTCT+b6xnqEIC2G0C0Bky9hHybXOuObkZsXkdClZ0FTJ2oq
+8RuYN9YtnnmylUT/KQ2WD8Q5kTLAzqcQqvgcV5I4d7g8k5btscufAX2HtlZ/q5ztfYxCEC09y7E
NudFEweaPPsYdricZhS7GaLEKeO8esgUO7lFYOe6TkWzh9HB9FR35UdUSAT8hIxj8/AeWDoDKbjA
ompwxHl5ZDCeU/W2Z37xgmNcEvRQk2xCYX2qGJNFzhyA/co1RdzbZ1IpmVEUDTwKqdXwYRGrYg7P
k/7f36BLsS+9fMACUdj4TPJVmjtW0ZgTKbmyiH/u6E+MDRW6D7GvtT/t7faHqZ+kZt6tZCCFJI26
6gB6FvaOUdOC3IeWSjZdrxZ3hnB+B8wXs6P3BHksXlLDRumh7G/ps4ucxWVPKmp9ijNGrjjqlN3Y
Ej8mfV+UgkwhpXohYlgEQ9Y4rjJOjaRL1IZtCRSu7t5/Dzn+EqIOY+eX9veKfl43OWD8rY/4Gx4Z
SPw87sLUMN/0+IVMg445/m0Yaq7b2D0UUOyuUw7ZjckYKSVtxbgWxoCY8KrjqIr1CETdRY+j1NbH
goqtpiEQ20vLhJ0RO0Nn+1JvWY+AHaQ4X6D7EAXiIukj8zk2MRtl+huC6Dyxml+1XWfdOSVxGoJo
w3nP3BASnL/yn+HVCR9Obh6MyekuIRLhskV7pnDrA67Oz3k9+TC0UM1gQaalj9zf+2AmdmmgytkJ
BAZ+FRo8G//iulFQ2rE34Uf/eIGaXjEwGuaNL16Bo0XivoLV3cMCtSTnh32iAVClBSZMOVIGgL5t
Se5ucnNSOh8qN3OJ1VmJE9qYfyMHyhqBZcZOdhf3urWHJUvKBGhFdka4DCvYnzxX2YWAxflel5MX
QmKPIqxCI0tfipDZyYDR79iFlyLOWDilSR4dRbWMssQyKMjSDBYl14BHi8TdSahqH6xAYYXrTQ+D
97WhLmj8x9g+amSuXxKZYo8q6TifsoeDv7W9sH+QBnrZejkUfEsUj9qQIPHJf80h5LsKOmCUUbvd
MgY6VIn0mhvEHebolwZJ8QaqM0w46pPnbG70M1Q13L42uirt79emWqzBQg5rX968HhRzoN25woXk
KpC+R07MFmwXBJDakUWKma0hDgarX3tdCGHSva/N7Z1yDNXKwpugX7aTLXcb5HNJiqOlrwJprxAN
OVDGPDY40MAVn4L+ibv5XrCndlOhWWz1/skuIrIjueG4YgEYKcluZrGHCASG/4uaR4Jnu5k9XrJN
581vgWnqgxK7l9lSkE18Mf3wleVtwxhBl31iWHBll/ms7W6iq566k68pVExDg6ADQDvBiO0HWK0G
EsjZo61K3kclSBB1NmZ4ADcUYsYLFPiERSglDuLbJPDK+Brm4Br8oA6lgop2hrCy6FhVUaXrKYUO
QppI5ytEiPDVfCJGmGMfZzFj1kJWAIhLOWPNeytioT6gP4amSI9WtiHES0/yYQYWq1M6KGOIHtGx
kh/5hzDIxIpZNsBUJ1fRN96dTOEnCVEZquiR46XRp7lydtnF3JXQrptbGj71Gslg3zXTJCAlcLDE
BuNOcGR/19kJWTJv5aRDY4naI54SkSC/A3V0Tro95Gp1OURzJt/Hpa0/vZDgAh57k7X8yEjnmO4O
ZI72eDdSLh6pCcFoVMYxzUv1sv1UZed6Of8yUWvfLPeivhrYiUDtXfRs1s+NPDV/X4WJ6U4p3WUe
RzQcHs/A3N4LVCZFHK8Z2SLeJwKAnUV8ruo7yj7wCxjjttb4Va629MkcY8KdK95YQGIlhFlWlNaI
9BlgClUDGOUi+OYGiZLY3cuh/CjHb5WO47/DTSiBp3a4kV3gczo1fPdu91GPWZ12Ut8axXuEk+9p
X2QqXbUiMVbL5G4CckJ+Enr0tGB8Fk0sUms/2HN+4x5tEHZQ61PJRSaAhGCK41eX1for2m5foXzX
ImHLdqljbM7e/KcnZ0x/U6fNpMmJgQTEWd0jZdmUyBOKMdYqjhKlRZTBrTPwPqVY0zA/B6y3+/pt
DRi04k+H/PDnkVMUUvR9B1Kvt5NCO/wjrYuDPm3ZCQXpHQj6AdQJcagF1TLHsDqwDPHOdVZKJxwt
NcXkVCDwi1vxwpfk55HTzSZRFLQ9Op+OPTYVQmbn6rJ+GwdvpQC6OMubNbRfabGK8mJA4asmSuK5
5s4NWA8PzbJG3WwkIRh7PlXLvgvu60n1zjlznhLgyKyy8okOwklrpH9vZBe4tNGTZNjDznCfBhlv
akIhrioR6AEcivnCPKqrQ7SRg8zEhX7ihonYMz7pbe1tX0Z8BSl60/uGDz1/uNegFuDt2AddRC3y
0spc47UrD/zg0s3PcoCYecKnNXRyVNSRW5gfsAS+Kjj981g55QyYFJ0BbYu+vO1JPe+pFVtaFO/6
c1Dg2/A/JCVhUXzGlXFjMV0NruW5Hb06cnzFkzVtkz+p/7bYVrK4fv+QTMsIBXtSLLogqJwIn7Jb
90jJuSiO0CgJzQeQXcHgh1n3IJz2CtptNPKlAuZUUSnb+9KVbAEkTuY3LkXWCnCj8+6/mnxFZsNZ
LmsfuFtBkLC1eTD5cgUzgpMFOnsTxbV9KhqocWJutwSPgGUGPNY3AQElNVRkpG2MSSK8ffwRY8n8
8vXWIG6e+GMb27dsEaG+wEc+CR0NcQCCmWaCz3vvlfzAb5ph+J9zoPxH7ZcgbR9geieLYrhrhWL3
JJRAiDLqxNdxk0LcxdcoHNs4MX3eo7QCYKe+OQTGcWgE2ojjbF9H4oBKm09yxhmHxwzvpwiC0phX
cPFgiqXbc16RXgSit+p2u2Ad+kubQWb1xK2rhcpykqxFvXDv2mvZ2TtCebqj8nTGkK9U9XL/MVkE
1nPlvDobS1eU33ZWtjStAsz6ouD8lLa/PI9qvO4ZPb954Ke7B3j+GyVKQa2UN8uaQgQF5PuNLnQW
phh9GkQ5gDr9AO/PZ3/e/jOQc7z8VxRdcKxYg0ckCE5UjpJC2kZu2NDtHlUQKu1jLvS9fk5w+n6V
jKq1jmyDu0thpcPggJ94jPjMnAh2omkTP4Obsh5ksQwTDrH0RHslhSGNC/Ek7PkQClA4jCPRDVux
WX7RnUzrKETPmDvDm7LRmUvLm6A9UP8uLdfM0VkZRiN8EN4zd7OubDFP9nuwqQsMsPJXS2nK+hAR
XwBaYtzS63PBUrS9CL65yhvduCNJn/uiLZ1qrklCp14LX+BYTa5qmqfTFpaj8x5j+AiMDSCxjjSE
TtqXiVDMA8Nb0S99sZxO5TgKImDiFBGwKvOR/mUk1bFOAtamH/647L5RrCR+xOF/2S6lbjG5OdNY
SkkkTEJgX7Nqi8twqUmf9vO/4Wtlp/xvhAVigodPNCU7Jp+gxpc8Pt5SDY8VmARuNjsqCglC8g3y
2zAFgrgmwmvSq1JsZtWXveYUHDWqOq/PbWZN96ilfQAuWYEmq4IXdvj+93zMbSb+RVWmWqLagzGB
rIrBwA99r/Mehd3o0akHU3vtHS4GNYIyKoZbNaETH/8LfECDkSs3EyFTPq1CFT2lnG0HLkBUx8Uj
jhSUQYSDaa4XWRAHSRosldFnnsM9b9kxkbjrMpKBJy+LA0F5XY9jSwgIQHteps1sIUS6nAuOrVJY
Nbaczse8FnKy9OdRhnq5kJYyg8QQdvkyaDm9VOTXGuy9DpE/lYtZB+E9o8JHyE+6Bdh2iufqSGNo
4wcyURMClIQnyWA9s7OyqbMvbiCUYxyw+UGHZMsKPLjY40+xHQvM0Lqhc4INujBRKv6pgfTNGivq
z5rKQcWhgSkTfLdxgD9SwsluKZw4hJlf9bJrj5/kybEYAmXxAWvM+a0lzFk53izr6RvaMl9AYgvU
rAEfV3c9F6KI2ke4mTaAFBMUpAsx+Z+J+BSu6J0mxhAkWRrt+5KuPkXe6GAT29NWfbxiYJN30e9m
Gw8YNAffG2XeS7hnnm7EUvaeDAz5OtHCVSIStElE7Jz6X8YkAIsOLaasT+2HAZ7jP3/ZmF+lRdrS
UTGoR29WSOAQ+bxWE1QxUhlKo+4HMIGZuGwdwU+3+TewLFLfHFSrdnvypnEnXgpzmJAknda8sXCR
GPHt9yhvXdtb4iknOCogk0cAHXoGfHhwGMjJOxg/i4cK00wRSkMxE5uxe2UBGRg1Ak9J40Z0E9WA
rNx/h/oeGgylbbxiXz/BJ8SgnPA0+puV2Nq0vA/OkPUuq6G2cG2I80gw7SsDDRxwqf9FJFO8ulZ1
4TqFGVV2ky7Kil5ksGGImz87KD47Pp3d9boDb2I9eNPELxOayrL5hN9wcPkL6MmPUqj9XYmeaQXG
ag2wLeEpkoXYn6eGwxZTdg6fk5IzrbAkWlwaQvy+PQD5eWDpq5WWL34pFkpAmW+c+HIXrsf9/Y6n
yeB6WwOhv6QVAkYAD4E0UsiDsjOkCW2HTnmzVEFyGKkbZuUcKtUA5TSNVAnV0ph+1umeCphL6lK7
0ex9KbVZH3eUJEDuVlAE1FRNpv3ZQYg4FCdBfz3xFHtgwCg/eB6PaD0hhAoGCydzaMTyE4JZ+BOW
ifwWKCmI1zrn5nyFz0nuLIuuVPfLVn7Dw/mSxAhLsiXiWaE/nQzP14MWggBTj/2tzEqyGksBOZ7/
gkMfjx1Qktq3fUgsk3peC9QNV7Dm9IvFGEYOdYfYDwUFqgmR55Axl6Zv5n6zydZoDWbaf70LLvV2
38LVti8v4dlCeORZ6AZib2HPL8f2d6BRXnAsdnhuKPCAhp/RPbqInaTSAnLBuuus6B4Jlr7XbvDf
aQCgm4ncDJL76f8kAKwQZHitUhtQnQrL1yYUDeE0HpMkT11Lvr9f4CSVM9BP/CnaAidKnhLlM7PS
R/ZjugYT8XegFo0Vgi3Ka58lH1CvexeC+IOudcwnNzE+tFM+u8KmIDLOZKlO1zN2QCy8II5iAzSW
1IOYOpYUTFbpfA05B+UuLpnc82ZBLDhdqRd0Bzxur8BLs/j7pvxp6f4xb94JlwjlM0ItVgahQF4v
7QL0hzdvWD4lyIQ3HI8DaK0mcfDbdWAt/nFUpZaDpVx5Q+hVFoX6ythU0+m5IIehkpsYgjMgYiLP
XvuH93JeVFi3q0mjy8Hm3IG2dZkvEcYNYY13Xv9uGlxfY6zsz3V0qz6LHhKpX66AWgLwec3fVQF4
DZA/7+efa9GURdz2iTxnqvQ8cnZASXVAddM7M6W7nTHgFvSBj0Gc6fcjdmUcBIpdOJO9+j4Ebecl
rY0zH/5UCP1+OLCDv1fb47GQU81SG16YuqH0gJ2VPlQ0snA9uCwWH1bb1ansaqVzqMj2v+qUrnY7
IgJ5S6hfM7HwzXP0lCwvJJCBA6hMNRr6ydQTl/24aJZmqNWdNCUGl3nMj0LMoiJ5i5mcu79O6F4V
JHjELAwtr+JQhBtnkC9JVbojwliI276KQW58TlMAWoJRHCO5WxO2sL/7TvXVoK1moSx/Eaw0Rysi
ZvPkZ59GBpn1WyiglYNNlCbA7GkP2f9QbHbSdRIFV4fcVNghPNiep8MFZO7Ux7UJghMP+9nrNooc
qNKFSFzVGbKGat+llcW06QUwT2e84ubzkbX0KICF/T+ELjzRxjiFzw+J0oW/hhauE0I4clkg1tX0
Dr0RuERFCEnhSwJtfhpvgQfO1gCMc0mvTAGwnhhZocaNo0jzP0yegfl3VZ1+EQPelc4/AbR+1rT3
ptsTNJ7h289kFdsvx+aQyD9aFcAtkhBY8F2IG4t6ht/Va5A9MUg1JtCEuAWb83ImDXy4yAMSxrZS
qUeuruHNShN7VmSoHIIbimW1O/SHWTm8MkjKUyks5mUqE7M4+BLuS94jQCdnwvF9jdLxSOPC2ASi
mJhND36neDINqECbAtn8Qxf4qoZ05Q/jC9jXcfvgpW9I/pjdE4v3PZYo/83tTjPbzhZ5u0Fsv6EV
L6JN8xLBktHdRR/bRymjmJzjw1nKVuzDKDhcPmbqSfU9VYl23gj5oDyjjshnBWsB9yYvQ8TCO9hr
+rlfvZT9BYmDn6rLFncMNgNyVSiOPFHnf88QTYggvuCLEX3Ey6E7TUYG0O0VPuAPNo+wV7TWylo3
IWiDgpUuzezSgasGfxcMzpYOPOFoqcrhOYI2PPfVz1zO78V9FNfhcCd2xEKYCtjs7RNCHygYRell
zqp9+SAr6qx9wmhzHQwx+km9tlaovMsuXkolcyWqzEeeqtAsoUDDX3wKI41zzEq9LvJwqOFsax3u
LVpWAS6RaBjA5OTjsvma57pVNNLW5cltY1sToZW7lq5UM22cNOW4olmOu4oBITdFVJGCaX4RykCe
mBM3zZ9mlLGNHYZ2aW3ueZ+PdexSBJKti3C/+O7+t88oTxhSIaOPC36T+PjFLveKxPPoIPcKgYyV
ta3cCC1jrgfz1PxEzK1oLZZKCPjr0/7AduVK0G3rJ69lmcsCZ7E2oKrLLIzwTjOvNK4JJhBez7Hm
uYoRjIzVtkLiL/1eu/qY2v4G3y56rUpqCxteWiaTpQyeRuXWwdHnH8MGLweHNJz+Op4a3FZMSWfB
/dH9Mu5lOECJU7IRQgz+H0ZPRe0PYgdkAXvsQeZrkHhno/Q+hRtKC/X9HdGsnT2EJ+Bi1CpLAa/t
XELzT9VjuEAg0SdzyimZMqN4KaHgcK9+eVQPrJvEGmzVW+5OKJkaIEKw0o5u3rkUzRUuGJfw0gvM
fo5CX3Um1BWc97Y7wRNGvffCDirmovg10XI7jAJydiMkSEv/skYpm5YBTA5YIffcS9S/bPYIcomo
/t+dExofloDfG8h1B7Ds1p0tpS+s5sTZc+0WpQstD8/PQURwJG7ds9VguCA8Q3rnui37YoSfhTAe
ZPNx9QecVRF3BG/UUrzXgYLfrL2mSlLbY4aO57YPukbegdNYlZcbGfN3YLIOZAdIqTLvGNy7oYXv
kvS2WcbUNFxMHFdrtZNkQH+h1jesEdvtktrUcvipqZBCr2U0+z1mhkNIrvOoGdm4ssjyqXJ7mVl9
SoOddWjoKI3MiNc2vJcMW3yqpokOXcPLHn6rH6OJJmsBry70NSZNz17dxEMyzbWfoN9FMveZ0f1j
H3/dDXkbp+tStQ9ifPt/hxEGUKBq0n8b0Ui+uPS2hCZmdU7+bHKBBgQRXtFo7AwKoh1vH4SIDRam
7J6bkNUrHNnMo+Y0ZRwUkQngPv9Sel+0Iw1JwOkbZRgdrCp5I0Z2cWSFaK5aDpHrcOxC9soMAeD0
u78yB4SYGkxj45mkSpmiyvp4Eo9CmCNjz7zl+kWrB3L9y2Xs3T3m5zD+V1vgIxjXtMaQ/sfjm1R3
mpiwhllMYvEgfCWaFfwkc7km9vPytx2xFWasRkQUJN8+g5C/HGYIoBPFu0S0mGf/185f6gPOJ9Yv
wJYGm75ekClrWYpFZ+NM8Ts17xPO0Ao+lkZDoULMdfDmDbFzcAxf4/n8k9Oij+dEjAHltMEnLHir
MWir2OaZ55XPHAqrrotshdFknZOMFkobq5QUxUSd5ImleTaKURPq7G2r5VxLfDW9uwvRMHLxRFoU
EIJziPA4FV16OQmagyDBFAw9pjyFis37tOdVpOxUJDS4BTcgAOx5DmW7HAbOCWzskHsiO2fM538Q
jrPQq6RD9xQDwEShJMTYMZnxw6lgb+AnHU0ebjdeVePIcQw9XAGbz9Zao4M9NvGvOmJflopy80mJ
c2KyI56GBx1jRdIIBn1YGM2iOPZTWdj9Rybw6t1XvMQzRbeEyaRVDDJwu/GBwKymK0AT+dTJD9MY
f8e5nBPMZvlt+JcaHTkpUA9SMf6mIGbbaG5QhBm1j6QlFFaB71KQ5f+Lv5MORYGpBi/OVB+2fFGw
OxkDrN+elNohGueEo6y7UsU2fG6T2YeLEiySgzH6TNViQVHnufrZHyuNHsvUcn5vdr7ZBjlRiEDq
OB/ogr2T2Dcxwjp2W+o7UlLnp3JvNKciQ33dW4cDAyuYPGgrhDZ60Kq8g9LH+viVKsZrXvAgCSKR
hjMOXxd3scd+uFMeInb4M5FrXUj8epa3HxMud4Lbqgi/En7AalmVrvRyxqJOG3mAYxOga/VNkQ8S
uTN04DfEaKpTHZA35gOb/FZ0TSfQdYivrpsXsLxWiLSGV+BjYTCaRTVX40uGXALc7+wXbJdJqIuK
QAoGzIHgCQCNv/tfkW01ZG4XLB7rj/BpShaE/h1UbgtXVCYNud/SuXPURN9yo3oZP12VXeevep9a
CG/GIhDEKyyAxDan5vcOSwNbzouz5TmJ+iTyZRT3zRn1C04nUFutkyFqzT604lhMExk8QvMkfAGZ
7Fh8KVMIsgE93mQl/S+MdtqaR6JtyElesnfSALM73PSkjoYHAl7TzES5MoRmOjfBqewqhFwYynSV
niv/0eB3aCdiRq7A8iXDH1OZO8lH0xLRVdnQ7xc/6YT25BC9EBSo1nCVRVL7EkIzXMO15zXgiJBN
VtS8viJz74zIXDN25qZInqMSMYGcxYpQstaBeEIuCgnznHKAf1zOd8iuGzKpBm6jKiIqTo+ccIpr
k3KzbWOcv0mOiEtRPAjnw2y7vqFKGjyhyb0UFjOGpAlKDVvWyLqmwYZS7oADB0vaOs463P6Iy46o
J9oO7eP91JNtGkCZK/biXddlHpz35vtDyixlCUES8jeGZ/q+oBORmaLmf/w9Ys2Mn+q0JbFDnu0e
oIzPLCYUkU7QwfmBVoGCHg+QgNwInh0/dl9Th9k5pereplieC3NN6M+sg4i30R6RjaMbg6WYNQ7b
Oj9SNL7JXjuaUBCzU7IuWczAVRth71GbNdiS1jdi2Tad4yZ9rBPevXtdPOiNrGapIvG2eEd9Qj0n
d82ex0G22Ulpowtc8e13SWw/0a9c+K91/QN4xLBLutGfslmXqwwf1baA5F6EoPPycIUWjDlFXY0U
Pwrw+qZ2FoE/IPTm2h/uld/hjd69yOfY2E8UsN1wCpJcykFiQpx5LRJFVoc8/JvRs6EkR5QBc1SZ
xXneyFUsZymDPPrdRSmKIVE9JU2iuYhFKhbVS9Q2s0BNbvojPQS3hmoxTmzz+FXOnfNNCxxNjW6i
IT3AFVjf1OWVA6dpDkvABFbX+5y3YgaEzhyDEivDxs8WxvbUdBSYLeAjXBxnmoPWkqJxxFRByOoF
XX2J7g4Bz9+7pV3M9PT/7Y29Hm5MExr9b80Ptr8Rl9n6yrmrfmxVws3xZtkS32zG4cqdhn81suE6
lk9vcHHC8l+II5D1PH24cazAxTCI1uP+1MQOXwGo3qJ+qTzl9m+/qpP0YkJR8ylFYju4FZhaTcxA
94mMHZfp310o4A/ldl9u2wvwerLX3pHhL9NPApKKKBB3KmTYra+8wrGFvPY5uIbshVofepGd7+CA
U6fGA29+MneK+Ls0LbChrpHez5qquPrchbGY8tHCm81cBQY7xlVbuzIGe6L2l+EWl8cBDmwpBBOO
29VJUzo+QfnlfY3Dz3eP47h7hZ4ldu8XMhPGxccO4bbIftJDImLpmXXpxqwB98NTdtSnvKzsDUK0
wa17X9IQPPE4v/Hsy0hncItk5da7c83T0YRflhF9+MiQS52pCFrgHhKJsVmcRFze5FnaY28Stnhv
OBQTGkAZTMYMD9SpVccNb31OZ1QF29n8kgX1bhncsrrYcuWgJFQosZhvMvLOl+abGlxubTrBUQkt
k7BgD4X9ne5VVWxZNUmNWGbZMbf+j4gKQY95xY27ugWNrVhFtBsvST0xiZm/j42cAhkn/d7ULr5I
pKpLhUa1RyulHpwlRzh7TeBfL0bVYsMT8k5CrQWXxdnqNrjMyLdp8uzJpWbvtJYqdA7xhCsyYRPN
poTI/8hUjNtnagIXfBJIzMmEW/4qNLYlHWOo6RvrTirmBpaqBmhsUINsMG3sIxOxV6fy1Oo4r3GP
VApJwOqiQwAsjF7888pZnKM3B197k9vGyJDkqdIQuyyK2j0ak7fBEZp9of0AQNYeTYfsO3uzwQE8
bV29J0hqABeIVmNsTAqCxmNspypt4/MrsrzrCMvBITMYqorCtezXSgxg+lYsLHmuSTtvzadxkxIW
SUKQIfkwvthYZYFNAav9/1jyfCZpNjMdnOghbamvGwqZA2by3lbqOflw8pZpti/zG6c8g5v2ut9Z
2vwY+KwTG3kZC45UxM9y2wfwfZWaPljsH2vNsThVb34Sasf5TjHjYIxDkF4qJfVYtnNI+koTF7+m
jVq+xXdEStjYFuZQmmL/bt/1K+rgfy/4URmYkuglVBSR3mwhWJX9lEOzuCnRRhq9JnvEadYDU6sL
Tde69r2sbzVuAH+D+1KjgcoyijYlpdkaZ9934Uh6y4ikL0NT8fcz+6TU0Sw6nvd6O1ZxnsiCcpSm
M6kbdBJFdq+dXZlxUwg/70AMV4ILx74RshndoSqXPhSkogSSnixoikWhgAmcPWHiqgRZXMQgRMy8
WfcmuBvIt7BN/tKdzTexwFul6OR7nl6yD20iN3EAJyZYhuvr2mJhOexVUiGl7zlO738duqsnFq/m
4x4lVL0aJ0lvXB85FtdmsP9zIg4xnAsrujoQY/BP9b6VxdiOOq13DXSM8GRZQT++itBRZ49PTxw+
wl9LmKofPC9UH1VSmR70KCZXVVtBvrm2nF7XVT8HapWL3buRU5Xp6qXJVIooVhxoFZYHNr+IqQlC
tCbhO6BxO+BOPYUjmgtlPUBsXQ660oxPzCBcupXxOcbIfatIh+t9Iy5nKwP2F879xvpp1zArYiZD
u85SYGXkf1erdfQzgljdp3trmU1q4CMVT2tEImWbhNHRGkEueNZ2pC8Q/SZvs29m45d22t0JtXxc
e+VfjvEPtB4uj2eYM5Xv1zFbkFyPhaOb5OTjADxBcOBt5NuFyFDEMoqwM+801h45f94aJIh6xhCN
fsqy5tklg6rKDzDAn5jyZsVkHLBABCZOg0okCUOph8TwEfVyT6l8nALlAhPFn4hRmpe0ieFWLn3V
Q8rZkKF33Y61nq8xl7aZvToQZ6D04I6aL8l8hkEOZd7uQ+5X313GbhnNamtnLT0TPgcJ/6u6PtMP
i8k36+U3N7J0dX74d8yw93N9qjuhdkrKJAiv5QDsX3a7GmF+pMaTrnVkM/yaKyVbwE2SbBbbE0jI
BZfG4jXJ+zZ+jcV+ZMQ0S/8+RdidyMyMwGFYnz5iq1oktIit0zLbIAkuLuVDuupWxIO7VPOA6Srl
sNQxWbrum+7ZrLMsD0qKNRV4fcAydo11utNxI/GlZyGbKkycO35LCgOL+3iSXKdjftOyOAQgdpk4
NgR8kFWTN//l38IePVhuY12yDrAEoLrcq5DggPXde7DuTrYXhSzcl38XxfaDzqSRQdc5p0ZiyK7q
VZ6oviWgG54DPg5QlRUHQq5bxZCSGZgtnJJVMKDJFxJkEmETUJ9Njb9AcN+ME+KUejScgvQx0O1C
1M7Lc3PdEKbIfre+f8f8hrQDwyVvpuSZbfy5tkBeboZCDwzOdeBRqqxZnrpqgAX2/U8gmuLgFWCc
xZkKm8yOmJST4S0d2DTfxjEARq+KvVBsDC7WK1PxmN/4PlVI7FZAeFU3QUs9uOjtac61k7tDEuDz
/XYv+g5WEi7C8BB3SEPg4K1H6MT0X2r+wsdZ1DZt27l22Czr9fUQLpb5SOXRV3wyc7PVPMtgGKND
vKVuHUx7+W8ZgROwDW3ChDi+yipWDWiOdu+G0DWojb64u+cFTDdcC7OTEBBMfSD2bysKlmT66jjD
YClxbKMG2qWiq+4WiilDzO4dmO4moPJqPPI6obuwOJ5jHm93F8ZhQ1iC9pb78+qm8Eqrsv5amlcH
k4MM4+2KaxyO1S4E7D6QeDXGFF/QAciB/KTk6x2jQ+JBcUYLEP8W+jm5w41w43dWYnXpirOucioB
Qd6UdpImiEoRLvR6Ya9FfJkQKwXQ5J+McEKaKddeDaHU3FhMRKM5XynPwM7ZYzZfbppuAHquqmPf
LJygwoEtOIv3C6czJ0K4txubLnDjnIWjAfWbS9ySbHkCIxcKllSO8aP3rI914402/VktmUOXKYkT
MF6uLxp9OAcV9r/8cCwdi+PfNCQJszmG2cx1ckyj/z21301UXOUnWHmIC2af8LyetfKv/3EN0FUK
N8yD6xiwi3qt1ZV04e5FL/pkm0G46SbCZ0jk4rsCKXY+z6a6bxkiyvhNzTlTfbD6yBWRipqRSt9Q
GY9X9gYi176BBVZDQtr0E5PVoSTws5xNvJ7/9S48aZPacIyQJn9Fb3rs+gfJu6SYWhBQ7cMUSDgw
tb//cxfWwW+Cm4wRAVnvqarGc21647rJXaT55ydomCfi5FJCvG8jtug+srH0DAD3tqo0pOkenM4K
fz0pHXamB98kQ2+gw8InMRVQDKGXnd3g/oOOnQqQE/yghS1uy2KwqetVn41x0viXRzc/6hWULJYW
aqSB+FEi6bZFskQjJsgbL4F7vZBHYzOQEe+yrqlD5a1CdrtfSZXF0zToVbqL+amnG6QfwW2BDSG9
5OJxZMyVSIlwfC5iETrpj2j0Dn2yDQBaf2cZ8XET3VWMWKx9ffDA2HfZzk5oS/ZoINlkl39zKhWA
j3nraHZF5/8gNtxNMRDcKxyfIgJS/IgEGVwPtVnQCNLpjyv0hWsGDYBuHbrIEdE5EKi0MEGKqWXW
01mq+Nt1MjyvUepumj4n7I+n4XfQ7qVoUTwNcaMkup26ez2uVmexMJdOU0X1xJpzxnE7YwgFeH05
4U9DXfmFCinnI8dv9SzaNhrTGNQwstCF98ahW5obHgT8KHpr5p26YGcLfqtfmkgTlSsgbKhPy88i
2uBSyGVgjXZtfKI7+ioI9Z6sfDzH5WJY7DUv2Zf2ZlQSrf6Jw3hqrYhCG+0mqQR0i2LR0DHwl6xx
RWG5M6EVbdIL/m4C07hdZWbAiECeyWsGDOwuDpY08wCTqjYTEXuvaS3qVFtGqZk/TN3GXpcDns0T
j5A+UBK27ma+81JrBw6IevjcC2mvE++2uXiPUheLz89XUlJo5ipkUzfR1ai0YLKoTSBiaiiXqMli
6wse4nKFyhJ+94fBUU5nJfIYatQOvLWXjqUt/KMJNQHemiDlZqs8C067ZoO/LJpYtAzk3muaZngP
2nXWc3vLXgrvfHL5ZXROF3gqpwPLhfntW6H4OlRTGLGMreXdmhCukJG7Ygc2x9wmlsM1xHRi7eEh
tRlEQuuBJo2Kf8iK4WHpPKY6vFtC9Lz1SHkWgBRjf4lqDgPZNzzaITwNXCxtnmeZO0Zyk3x4A6uB
NHS5lxkZ+rdpBhvLjuydIVQIndGmHaGf9LhAQhDe+3Q2dggHTnuG8N+kh+dqkq1in6TAMYmfF4O9
9sdYhoFiFQU6sxoH42j+VxKwNeT212uae5U9D5aT7lue5BAJ7BdfAuWUJbU6AW8y1BJw04bWrVkE
II20ZDizxVGgNJJ3UV54Nzep+zAWAPaJii/KGudFENcjI/d/xgzgdBRghRE7A4EYotGuEbyTqrvq
FqGvN+7Ki0/BdHRceK+zHAFKw0oKM+HfQhgCJiB1TGXpP7aM1nKBjHaZY/gcoEJ1C2AZJkxWIJNn
26xD0+bxb+pMR8CYniFPIlNwfJYHVmHU59cAgUKhAY49KA/twB+7W5uxA+ucAzc4SfDi3qedgXQF
rYEpXmhziqtnfyX3Q91J2uQF/bMuupzDJehVskLiW8ibcaDtHY3/tVZGMHRiCltQop2RPU1YT/c8
VGCVqbWNAMmzNtOs6w/KUoiSuxjOkSJrfyReLiSnAVJ2zO0PW2jF4BWGyrpUKBzD8ALELbInsEdP
nykNSYKd6TH+dNRpKJIrIIQM7nn2cID1wwydLaZbK2oJdzlyT0Ef8h9C/264B6i2+Z4nRgQfC3DK
OMonKHd9XzgtVq6XcQF2k18k/5DTFn6uqBkHIC4XTzt2xPvUS0k0z9zX8wq/5K417NWVOqQjZ7ZI
UEGmT3rEAZxLo2BZdBhF8R4O2Z7fequ+tkTZMUNJ0zA1ifbu1rtjfe+sSyoBmE+6jE+vP2Oox5ER
aGhYAHTRaM+4lXNiiZU/8A+aE1YyuEa+xBmjVw8757Wq5kyZ2UhnG0jrI+ct1KX8UiFXwKDQSJLf
AfJt17FPhd7Beosg/tKWdHm1onkG/UFRe6/RHbgZxDkWbIlNhvXZv9R48gd2hZIY9U5+WwxCesf+
C6KA8smBGBWRCy2K8+97ROyPUHOxE1aWXmWveaBzz32SnUV/iFk833FvmfxqHW05OAk53ngbh+P4
tmWgHtKuA/9klG5gcCE4V6Wrygqq8pHvVPGZdrOL3gYEpNfgrThp7McLdXZx/4r8tuoTjZZkUXFv
4mGx1Uz9fkp0l5KR//wgYC3vYoJit5py45szZeNm/sIAP77+q1J4LNSa6AvP+NWOX8qNO+r13Z+r
hSARxLVZrnIPU+KQrAJVMwC7OjptqbF4SoAx4zcpAZtOVuOfQLFEK3oYxWi50WldfXN0qZhFahla
i56O2EhFxFh7Y4eoKJnuWHh8SM5gKhegcrq2xzXXkguvqHTcA+Jz+rnlmD/rJ17KjBYdNFbFlker
l688V0qZRIkDi86ON628iGedSyopaZ07Cb4q+h5e0NAGFSw1jpFqHhRbTHBLx0gQXIi99/DuFk0S
MokrlI8HaHb4CVCemoGY6oxkHjMz3n8EnAKYBVFwlHyNpE0Nau25VJ8wEiMTSjOwovTs44rGlWDS
XCmRtebGQpSBaPO7gBtDAXT719JX6BKiKbtOOMrlKsSAZu03UklUsqo/4DU5mvFO5RYDuIwi9vZO
gQOf1+M8FlrjW0BPMyuHNgJeNkXkM3CRZQ/U3oFZbIHQ6jI6uAdULqgx2Pp1FexeBRTSVSlSyrr3
6ibp3wHAVznN0/aeY9R0vjFYGbbXi1C1nPtNDBFsqVsPRRHa+tWj610HBZrzcbJ//YNsBXZQrKNf
CW035Qjn20x4EiKQcWXi/xJZP3GcR/4J4j3SVjGWVumD5aCo86qEBI64Hc/04QkkjWCK9KPWiWA0
7dv9k2LlVTIdS/gJ/PlhLL+0GW1ypwYtq+gVMDRA71tM/Ftf5UVd0QH7ceuoOqMMxy/+9O8mEw8a
frdoI3Nea+g80TktgSICIEbGvNuZJE9DTzbRMfFdApHNrdUToyTcDo+o9fsbmyYLcH7X3Z1yX4P7
ROntcCYYckjAoPhzfDQkIYUSh9bBhS3jXLVJJsDu2EL5DwLNcA1MWG+ATAz0lCnJ5Zth+XbSanhB
W9tU8OO59hZUsYGJG0JF5qJbhuQ07rHDmywpQACoDEgteSNAfA3DTJYHsVUAmaTuqwSMmNBuhzZv
yVk2+ezm5cA+MvuJgYaw2bNU3LRmSxoM6uVJR+efte+OoMM3ClPLGUro15yXaItV5iA3XgJ41b4R
M5h4QK6k1QoGmt3bZluqPAqSdHdCps/DZmLOhvsjac+8IxT4egIL5Ivd2Si+eXczC9Kt4oCtM+hZ
KyryrcIGajITBpvAY7HDfB1ZVAf4pOMfXiciSnWPQmJpWMQr/TzLXdVGK6Nc/PwQ6ZaAuqTFolKz
zLNx/C+UoKwOwzHSa0dhfjrZwYeOQ+sfP4YWCutSU7oEeHj5j1zFxVQXRAvOGRUL6mtbtTz2hM9W
MJMvLOtK/eLFjSrpREvvliG6+9q7YG/uLjK2VtfdygmeEGkJriHxhOgGemOCnt8TfggBuklUDGBX
2mzm5FEIpEh/YXdBa4UTISeLB7dRty821ADrAuHzvYtdZ3KK7kmPCMHbBUzLrB8cCOmIbr3sJHOk
7s/1sRMmBLj+alyOq6LrzlIriD8YlQ2IRYtpkeh44i7Y4u3GXcw4HID12oh07OCEpw3ffsqqgA2D
mdvnsRnHc6lvLOWhnSIS8TNnoeQrS0NGJlmwi1nFBDXtPuBEH+mSBXzm6G/QjBgK+sUBCGflgLhC
/RZHeHfO9sMkk0AorFzRjPPXNzu/z7mSuA2SAWEN+3m6cO7BjQw0UwmFbVS1fErzs6bULYKW4jJJ
q4vHfRhEW0SrVObdRX2qDejl+Nu+7TFERpc32LgFMa2Lvxo19CJSYkB6A6HQUdzQeEPKqatJZN+Y
aZj0lIhJvb225KUGHcYH5szWJdSF175LtKt5+O8v49jBGVSGjYWOChLwd3NGqg+oiVCZAkZOgnuq
eb2A9xwVvgzjKm2eeAwxp0WHQM84q4Z+3Ggje6jPbfvwzZDMkyUeKWh3DFLMPnAtLZ6Qa+2KowY7
JfTWd+nuH4wKErbXx2YhafKq6u2CCb2G8tsfaHZyrrBPbR/zLkBLXLEuxYRXBPku30i1DDIgbfR9
NRm5UQYnUbxFgY8TRq/J7UaDi+GV3280eC5Ypn/7adSkbwlgLtrhyALssSWvzsChRuC/PD5iQ7ZP
ZtPRErzzMMUq8yMHzOMc08sfavWlUOxVkZMvUgCQ+yHvFHDbfusBcK5i6zW9nqUU8zBB/4Tgzeoa
c+6ksbA6nSSg+9aZvW1heKNVhSHpR1m4+UhkltnYq5BKWdl/DvimWtOohdeIIifSXqkuXBXEXh6U
HKLJxZSwbgtZOXeorcZxmlPqTFG76LwPkwlKxIYyyL26H6LJ8ZRPTS+YKgoIIM7DcuVUKvUmCkSb
ENZzAgKvpXz4xVi9jqmocfEwnkRIuZTJ6+4DCoorZG+r38bapgjU8XR/LgFpZOKzbTHRKcs+cTc5
h0cRcBNabx5ZIlKJl/0bPprEEp99UR1XcH2M61mjpvEuue4BCJqiAZihdBdi+gwO1q6jFj+47z7X
7jqrxOvPgXqX/U0+GP+rkRO3NP2RDRHA4TIDOcHkpRIIg3PQ9kHucIhNZqdu1igBpGVvC9lG1M9y
aiKBZJwtBFgAMFsu84g8Vr2vNqVT8TEFtU2LwnbOYl3TzNBcA971c25LDcYtK/Xy2eVx7dMfIUNn
ABUti84vBeoy7J9DoErqcOaS18T6huuLJt6wQf0npOyGUTdDl+lmN3BOYIQhESPR/dM1o4IU8mpg
WC051tJqIeUBlzQmoNoyDpN1fDDr9p6kDoFqG0DBy+GCO9ayCt0eR0LZ85bCVxHes7FGEy/tFe1M
Ja5ZudNaQmjg65HTh3u5CPE63lrRNvAuQr3YE460Yefcgw4DwaDLB4slvUdI+tRxhmbLH8mpfHUz
kIrX5CQhWTSnaXILS/9opko7dzxc95qhdevrUYeVSG88iqDzutFcU9IbeZFBBEy6A+F5YiMI74Dr
1Te0b2SXYtzJTUIPkiiQbm3zd0ywG6UI0BXvze0rQinGE7BRfrS5Bi7wYS9q6vnBdk3XreL788R6
g+AI9QJqalFKYBHPSkYDzWGdYf34qdHor3fp6disrJnhd37Xg0jaZ/R8yq2adbhcwxdDcaFCGaBM
A23njtvMYM8tmiI/Lv2QuHz6zP3JDchARmBs6RbC4/kJFO/NCPPrc9GgHPHKEwtPMi7Wf9db30cw
2oA6uHGGe0jj+WIcrx1lCrP7JnXEZiCIbxApM5QCVyB76fsy94wlPYfZKk4ThIjgd/2jSOgoBRT/
sfbLf/o1nl+RAYNG9QcYv5NMSykRgZAkIRgK30S42oUnVaRC/eOPyX3dUlBxICsCZ3JSo44qdmhf
VCMFaV/pScN8xMDdiyZepDjORlSEuj/R8+0z877Uulc+wJXvliWRGpnceSnVyD6mGfbtZns485t2
lbR/lX97jrNQl+sk0IKCf/CauuHDsfeWHhLbEk45mBSsedlFMfrDP0o69PKBM3fdncR2v20s8vrs
lnTzrI8SNBTX0DjV6YGVBZgWll9hpNowBnwSp0GypeEXsIsd2kyYIhS7J5+jz0tkhX1G2jmMoS4I
a9pCeRmsOnxiazW0vzkePK5MkFcnwWWWK13ph0ZvzLxOaU/OvS3sYjZ6rNyYc/mkYw9tCCJfYCjI
0BrAyu62bCySlJ/ah4Qsb0Sx2GF0ho3bIsmo0FMWv+nIlkqrsE18PpalPtGxbgGfnTrmaB53Mydz
TseQ3U8ImoHkvphdnyYiGPAv49tEI8VpViKBeF53GNtCFgv7FfFNBfm9vi1u0EpZ3xRfoBQxFdTF
UVLAC/cJiRA1QzNNWz851rVNFKbiqp5JYj1IMzyP43m8hD79GGD5znifRxf8rHlCbwxFgJ29zguG
mT7Mx+VL0BIRqp9rQM+dMa2vv5TtwGqkSNqHlYlzD4ycE105L7i4mSC3UtznAdUQc9ER/64x9QFi
ne7RH5xkBDlY0kKYMxnyeowL7WtNu5RbWRlSyoK/kH4y7KEWroGTUPQ5XqMiPdhhOgFzZgqnXDBE
oOQ5Aef8fLJjRO2BGAJaPaGYk6z+9gf+zXZ0TwBDPItIuSEJHeSGmw/rPoSRpnLwrikiS/eAyXZu
Hly1GjX5m6PH2wYZzLQ3m+8fvq7P3WOevcuY1930ChANeEEf3o8et//E2n27uBw0cSMyt/2HboQm
Z7gex3ZR0slsPpHGlsFtGqgZfF0GHR/6GI+EzU91CAzVGhAryGv/6SrNTn3r6UimX3PR2MGAy6Z6
EXfKTqUl72mH7ocqNh7s5JXBn4I3Jxvrb/GlfgE17V9MRcQ1vA3Z94cRnY1GlBBJ5ukBJQkjuHWa
N+SuBTRUNCY2w7iQBa9jB1OdQZOwcwrP11Pn+HgGC27Z4/oYGkUHALdwY66RaPVErpROkEEzwgSa
jsdUviNrwSLAPE6s6XNCvrI3r25wIJpNAaPusEtAw246w8agvq7VOVeD6h7LzgO1CNF/bfB8unaX
c8TJSgKawt3KuTpFtuhMj0VX3mqThFFugESnpRsJb9BCQskA5K8UWPJIxP9JXD1CM+RcjTHmD33q
JoOnfmGjORTihNhW7a+loIDA2iESIXSSkGH5vSjeVC7x5BEg0MnOOVXTKu7rtsaAau/neIz3Wm9d
P5eCgRTHNaM/pmhHn3+Fue3FqkGNiyjAuFwiHzZquOlGTkuIqOD6E8GToMU51s5osis5YF86sTLF
zXEFfDoNNp0ENeep4TypjUD/ppjufM2n4QEbUhc3AojmC5zKrl4BDyFZnc67aKB93YK2PCMTK5HO
9v9ZlvZkYLjFTwzX+dDFMNtQ4vuFE4LZ1GjfDoqXalJmPsWGyhPnCk+4bmVFfKBjXZMxzADkqRGb
thkDj3J++iYSwCmQzTvk2j7lNbvhSmdxnjgjwajtaVKRpifLmnoi9SbDL6aeYHnHzPYwnLDbKNfO
siHx4pvcZDfLygRyMn3LBNoPw2guROvtdaZ3CZ2JRBCDWQ63Sj/yQ/NEstXj72IYIFB4Kcodo4iD
LgmqScdzuO0E/C5ZmQ4h6S2/NBYxmhSnumaM3hjjXOWphDzAy1Kk4TSYbHTfaiiS90mKchM04YLu
dUNXweMmlJK7f16Hv5TgqNA9O4A1EpfmYZc+DilC+SpRmtpeQgXS/v0nbO1DA6OHrDhHn6nZ4AJN
zuenvqxWWYoqQkA+dAR1Yl6GJP84LSSzR2i3cXvVj99bVFTJBFJA7BvFVkIZl2kTzxjn1R/Ci1aX
E6nhyDU+W231w6wpavGd3/6e3eRvqV7jLRjZ46uuLz5keiBInHHjoTe2JRq2YZcE9IFrkeZ7QCLm
NKJlMXMoSiUS+l/WQiTjGxCsB6RetHrv+RJeXCvh9uXYkRbBjrQakGa8cfltUAyjcWy42cTSBiTp
UqflEMqkbCrNy8oLfNwgJsSgAxPLphmwULP0/dVEuXmpTyo+aeuVEl9j37VhUYUE7/D9ok19lWYd
6q6XD3fpaBvMiMeUoKr+1ME+q2bFVVKEIMfPmMGqx9/Fmatdv/8c5zR131pflvyOLfipgFeycV58
eanbEr3mq+5bCpvpKtcRtDdAAvQh34ME1eJulFQqNJRUT0WilTX/tSyWMOJDYxzYAN4j8guXQOrh
wcPPiOAFC0PJy0W95cFg/bBczf+lyHiavCBmfZlsR50dJNYeslmkBJSLUWMcTH+rvylAdTinSv24
D8+QFP8IcYot3koQgaq5nYeGQwqgAuBocUJT2u8pafylbpDv6HYZqd+cPHTWxHGufxcg2zQ9viE7
agZr7D2cPK8cdzTq6k075xcV3Srl1BHv7kxz9i7x103G3g8CQVeDGIMoYNgi+44vtQ9iOgULl2pV
2hA5tpbC1qDWcSvFS/QeeyC2bsgm6JczBfQr4AL/vJu9elTMJegCRNK1NFblJeb/qipJwSVsaEpw
cBgnO8JtOj2Zk5OLTWB6EDMBjCrtUDI1tPPmA7U9NhGD+ADs9RWcIvoJfJnuubSmbRBukXUlfLe/
3beqTkVfFUuj/wccL/UwmJxDw1wpKE7MFfXWN+bjE2TeWV0lDLq/1YkzWBEgGfKNp1gU2spT5XpH
ST+4EheQ5P93PrkgT1ZYzlcW80/QlZjzZihz3sC8mujoBJZp9rPRoxhVsO/TKGjT35Jr6OqMUH+b
9/EXDwXupEb2v8lhAyePN5gvh701q9lupYNHkOII0kGRt8ALuw9lmbCqKfnBt1pmEn6Id9Q9IlgT
+Eh0Dntvkqs4soodgLrkSI+wcKQ/vpaFMN6wUp/+4RiifNj77dW/Q08tYoMT3Wa0tk09t5pjvhYA
ejT96TivKFgHVPjUW1WsTSsw4yS/Tig9aI1fAKC0pSiZ4DUPEPlUC2s1eevRZdtIu6rGv61wGKuo
d8FEXhWuthYqbDyykTWi9IDXoZ/+62wvEQ4hXHcYB2ybKG8WbhIt0ajLoiDUF3Jp/QNqYWZ50AGA
7WjN5sNvNdhD58OSKhOnIzOBE+QIok5pd6E+WCXl6pd/jutQzbQI/oFBJauL6me+ZIifhkiXOtcU
hdUiiovbL+gOwf0eOazR5M9I7Ccs7cl4J44faytOfIegeObrnVA+saD2vxhiCyhpc2n3tbjk9y+Q
tAFSWebjmc37fek2KgMIlUUcPovdY+7wvblGDWfQkspErwwut5QdDUBEH7bHjEdpXNIgzw2IiIUN
jbZAedT4vWYuV2IxJkXXogYNJVoZmeVbVYk7aotoOPsGzxk93NojH/cInaTW+MAUZp8/ZqAM9KRU
pF0LvzmI/ZdOZXEtrcQN3Ezrt+2M/PrEr3oWiDxZvIG9rAYgGauYCtEZhaVl5zFcxkyQkq2fUxGO
yOzYKoArshmVLYxYP+dNEBa4eTQv37UBuOpFAx1Z43E5zrPeb4mcfODezbHOYxW7sOKxh2B16YOy
zF5g+ZhdhRcxv9CKvDPV+nKnD9cYKCflb4eUr9oufQAhzUjXI8zVziVIyNArdZ52y6VdEV+Sp1Lv
cgJ1H3zwRylrVd/SFNx+zHBvvsPhqpDjjrhS57rryzPHhZVZaOw9m6n9jvzUaI+Es86oRrYwG5UL
mRmJLBApqOW/sw3HbNJh5eDWUB67u1I5Ar7g0xujtx0GMwICqeM4NQcLrOZAZGQuLx07PDbTtZlt
VeiqT+OdfXEVHpyne2J76fKDL7xLd28Ox0iFMvt2Si6EcvPNFXlf0GNn6gqEK3aF5K2o2qUUUUBQ
KxzUkqw8jKbDgsPNi6wxwN7Dst9U4lKzyCrRKC6fMoOFqho7FJRMaDtDafyyJ/4MzGQ3QRvSYYSA
6kKtI3vNZbUMg22722mImUEpFUekOxUCKUURg9OjyOM7cTrX4f9GvDDtFWI9pnl10jt+jFuP6rZn
k7hqRkrX+JsxzIK2fYk4PaFJWTnrtZbnisf/mN/uGL/rptQGUZfbWTN1RkBsWTl5X+ARD+IYfINR
HCBUI0od95yfpe/X1rhw4uBxmvgp9Sp+G8cENyGpSrj4mS+hQMdNPpw48zc/qCwDYvt2Nkt0SyOL
zxmTSbmBLg7Mzzo3ds8x8fiz7lOH5kxCNNGTpC8bh78hgyB44hgEnSX22abNAHSEzTqixG2+9rXJ
WKNIhmBb9/bp3MPeuYvhl/L9wxfPL7T7gwS+EHy6KfR25b1rpWwgrRx8LfArtfDgGYY1E+SSZtMi
1iD40O5a+TTY3hJZ7HpYraB0XI1Q+jzxsd0n2e7EgwXdrXLE7HTmin53lWSjTkXWR0AqYn24CJSv
agjbUQ6jjivAdGPl33P4KvBjJfhWi7T00xb4IDsL+NhNM3m7IxLy/tgU7rBXnnINDMZxpgx3XGLY
aLZ9FmAAOq4vYIxkw9yDExL/EfuAUn9bvs5QokSi0ilZeF0RCARrz3m8udZVsxLR0mY2yDgokQZ2
CotunxQpMFVA7q+HbaRqVzUtIc0ZSAzm5OD9vON8BQsEVr3U8VFMOODi9juK7rWi/+ml5yvRpnlv
Fcxt4XDPX0Y/9bqv5NhoN0iIG+kUz6jSpjOLMPk1o4RdKwDjdLzR2Ii3w++LgpU82ERtd50IN6+I
1gVfCdy/ImN/5dSorCu2E7/UiKdBhtzILbazAW9+YBovZtCt1Scp795njHY4osN/p04ZL4A/98AK
eawOGc0iSnK7tk1r2qJUZpKR643JEdgK23UPa4l2Sf90B8jEfArsLbV3J9CIHLqZ7XdCVI2cabei
HE1jWa7fB/0MCM7mu/lgMSoFgeOsv5ydZwrhTTqr6GxhwtrFGdJ7Q+tUDas/dsONOBFZ9LCSZgSY
Df6AJ4BbUSAqQX4/9UShJ27X0TRGdAG9eahAnk19/nX1B4xKuOUJjLD8rebRCD8OGptAVdRwnST6
L61t3GFBFZaZiP+RzSK6VqwvwsB/U/mRYICZTEE6Dt71LszJMfQ01bNepjnA+a8vrGlvCXmianAK
5f5Kgba/QOOLYAA5pInOnOOmfGc012b0T3up5c6C9SZxHeM0f6ZIqDsGvQM8O5mnYwn9KgKSYnWs
4LbmOx58ufdQEjM4tR2GbosVp+uxwH46An1noX2azE52AeT2sXCFSumZjo6ufFhq+BPotidrW/FR
W8T9vLuvQqxTYqhy8Mjn8Z3NZMEPZoXVl73rVOU1gP7wqDTC8bswtdR8cwPm5jJUqjff4ipSOWnM
CkDvmeU1LweybGJPHoUBQjIlQxzAxZHE/dk5kafc1PmuEQkmz5x2yKZmD71GjuvBvy4TxCafq3cV
RTYEJjn2hG90sW0w8MeYKpkdikNLf4BhQ6exaGdfzOmn+9F9YBeVry6yLMcXgS9M/IGRTNI78ZLE
NLmB0HgFxKrRmLJB9MTnMUw5vCd5ccyiO7VWqULVrtrh+3t/YCR52ehTmS4tJjtuUjBZk+f0lDLT
Zb59bPsBvxrxBijd85D6MWbsZ7c6q+65F9MrgkqG3WSzmTyfzT2soZmdE4GBTABaDbiL+BTZQrpI
7qtDHswgQf7qXAdz6itqYTSwDPNEd811yZQZ0e9U8NyV54oPUyLJoOaTijbRHesl+39dMXnkCOBp
NPm5EkkBiwUROqsT7kyxMmoxgcDimCrN40fP1AaieYvrZfkBpnGjkL2O/Tp6WcI94hnZJXVeriWH
AAQ9LLn0SPL/Pf02B+ws7kqYbRjisaZ0I2dg7vmSshAY8nLXoYbWkgfkuqMS0qgvRERLgS12W0kk
MVwVnZJIIXmAaM0KQOBw8gNTO70D2o6je5gwf5rs7Ha2iwvqQ975MKY238wUQHbt7ROxHnMHpIja
LNrB+VsvGNIiMuhNve6SukoGIAdkVEQ7YT7fezQtPm2micthmFFXeMirUqW+94JRdRbPFLdFQOmf
FFwYsUU1VInhLEQdXTF5csUhqyhnNx2INXaSK3wXaM3Xt7Zc2CAclTnI7TpfyZBZAi0ikb+j8lmq
N64bryHp8xEwciBrA5CXMJ05ndLaU6o+aTs2iFCRLNG924QCWG1k5YjySQEKXaHmmNyyPxTIPwfp
1su8ZLP+LNoMFrHNFKu6w9AOSWVjehV4oG+C2M3oFLWZ+lJOWOcUr5Wfc+a9S3k/qco79OeQE1r7
15wz3KsfuGAH1rnC8aiDrewrq1kXA2p7qbfL2GF91+AThjV30HZlPKYrTFq5/pW7YrH0IISdwgBe
yWtbv7hTNU6i//kZgLHO73zp2rWtdXvRGV5gRmE0HXRTVqgqExiOOTsuCGTNwfURMD+2F6H/RPEn
kMgYrBurEbaozpVbj5pqrMyy7jBBPjtwE40e/6MaPsRcVdBK4gk1lmUmHBFsXdjChjRYubExKW49
SsZaQ7VjGdj5nSoc/2jSdm7RDVUkL4nxiBKbpvbpZAkqR7mH76+J210k0xAJOAGd60m4ypz7mqJt
6MHVcO1pXzn9UbFrNaxrb5rvXZeVZ1a91+/WjjfvwCeypcjCiHVM0UWZPg2QM9JOMZLa9cpxrZWe
IlE72XHLBcRhIR26Ip4ZenXoclo04cdvd2GI1qaGawBK9pbQrY96w9KAdPotZNHEI6YRnba9Iy4v
bfm5I1fydTJ00DP5L6Xs/9U7e/R3TqLi8wbvJ+ZRR7LCc4eVoAvypFJc06/DWO1pu5LXcne3MSKN
jRnLei10FGFas1aJ7T6JCCE1bvsSJ/uARfX/wua9UPju6wzVSla4SXbcawQ8pFM/SiIL0ct1CBG4
BnEfBwe6XbRdaGd7gA7oRZNfGAzPRHVjSgfWShRsLyCunI/WuFQmDga2wMGwGnCnBQcipvysORuq
z7rKGByhIjqtkHlynIGhSO5ekNTkYzf5s1gv+nk0SVVR5SanbNSWfJBb8+eN8vVVf4gT8y+76+Q/
m0Ks2+tV+Cs2GSUaHFdt09BUyCy6hRd8zm3A8TWGSxk5KCCattEbj5lGxgRr9LSckgMwG7G92xGK
qnewezuZeHY1hTQe8BVsplyUjsJUejWibOoDkDtaCZ3FLRusON0g4EurFqnZ0VCqoyo6n7CXO61I
wx8Y3yzWXr8ml/9pa0XUbxTLZO4fmVs4ZcyFbPT5PT6LIcP6c/7v743/+ZgyC48iMoWgnCBGwhTy
3Z7oFCrfugdMxx7wLZi6XtN3zwSyM3jMeo1AbA6KcHTdsWyE+BgfI88tY3tvMRMbpcqJosGIrAg3
W703IKwxUyrB7SMsOnyvcc4walA/arkHmAJVrbRo2n+TJITaCFeYgooxo5OI0EzGP2sDzKpoCKgz
S72s1CFb3dwhTPG8kXo85csSXdY621NWal1kZVdBrUrLwGbkLPPL6Th5IvlXDn5Zc9LSiOCiQtcC
JdewgdfQc/RLYinpYw+ZJg56JGDgJP47HvOXk1VH5E9bY6hv5vKlLQUZNH4LLLX1b+6QaQo1MYpz
fGFbC2up7NEwYV96nnZDAcI5R4ksR5uLAACz0dUA29HuMISfVKdk8ABorCiFXYbWoFLm8NtGiRRj
ZivxIfgFoETmVSh5eZ23C81iPDUCLvmq0MHMSU6GHWzEzyswYyF+f87alBQQOjvxKZqYxUx2M/XT
pGeiUEN3VTTNKvOT1BZ0UM78jUunp2tVtowdG5a93kBXSskzsw7bFTZKMn2WoVRUzcShYYR9tM+d
pwM+ATH/vMPy2+0i/mOBKoqWcQjE+iWOhJvqYac3mTVwzppKZV9Cq067bmTogOyQ+LJos1NH9B4e
7ozKnCyqbzt9Dng8h2NeOEjPSViUuo8VmX6b6o3RymNoYdKtzIC6z6vDrGJcvvlgut6vmRnlhOAs
BcIInQya4aQ5tpioXk+jaog9UrtW+WmKy4JZ2v3/Egxcio4ycFlvGEjkX4rYuXGdr82Wk6s7MsRG
k0HvbDaJH72Ls1XvKE1sSlN00t7lXon6HOhV/k2t5UvweRhfVbQB4CIWlcQBLnodL4vdVKphCXJ+
OOEmeXUjo6pqnLPjQ3Rt+O8cULen4AECpdPVqJ74VTPD9T17Og+1PfZEhli+OsWelqpGdj15E1Ww
v30R01dGiGcQzUasVjg/I0ngcSu8ug0BqtZyBrq3mFVwK7TBuIU15RPjHlHfawHRuksddPyWSC5B
8yTogPGAsFGRViXQ3vPKEhf1av47iC1abXHJ+tP9V6J3FahAyo4jR1uhKkn3bEH7n0Lxwkea1OaX
IqBj+BX5akAHHC8KVU6msLNYvjZpiNV1XzTYrYfyyhe42k6j38Galu2DXNMOfN6zZfcDrIevI4pJ
ij9AI54Q+wuEeDw4g9511mfWFvtpO2Scw2zMHkMJU6hwq+YHoNwMDhglysg7CuBoaDf8hvJfCne1
/yQ096vKUzIZ4OlFeEmMdEmvKG1ZykVr0+i2L1ffs7WlptdIq36ud5k995GUdo86QAFUQKnWEGIe
fXQhPml+TvaLyy3/jZLjdHlsD5LdQO2+3QsFrAKhJGvttlXh1o/I0QMJZd+JlqbSBV6xmG+ghRMQ
LRXEKg05EFjh/l9AK/NZRNPOWbfOO/z9oq9RB0s0LoEb8fyS4tEd01j3HmhQAXUhLXWqtJLLdWUM
Wbj6xg3KTe6KuBDOqRrdxTLeKR9aN8uQ9nkiYMCgpdwP5EosVme6XHhwXQvGUVARHVyDmPTtZaTT
m330QvIa+EBCaFj9BU9DC2jmX41XJTesb3bDHxhgPXaMbiqcZROL5N0s1eJ/l1HMvLVkyMqVhR2G
ASdGFXcwd6ygtkIf3cvUOs78Q3g4fcRLc+QQz5l1N2zvgiXnQiPBOZOqkaKYvMq4WkLD4rHkK0Oe
tSXuQmCYmVlOZvfZZ/PdpcrRUtQhWAY3Z22Nu7Nw2H/JsfPLlm9tXpiMoOVQjNEyF/8K9RWC0EYw
7V8mvQmuryrL6bA4eyMI6QqsgA7L5FQpPulxhyNx9J/wlvODDGVqGSyg0QTJ2keMINe4FwfiB0HE
pHUmnR1O9MhwVnWdtNGPETZVxe0IkzVG4a4tVCFNtTY3OCvE2PdRVIuogVPwVPHDw4XDgVGWzkC+
kbhvSvCqnmbCs+R0Wa9ytr+dtDD8IxFZ+asU8Y4SFWoY1PxbMz0Pu/LyibyK0/6w9DDaGxRySB/J
TM1W1ZN7Y+FFZ+myTdVwYHCkHUUiRW37dFPjNJRuL7MHTRseuF/nPZwCtvEkHwda7bq1EWCZC/sc
XgkC1iwl9+u5EgxCTYWn1nkkuymqnaECxp6CFVrATLp9coQHsyXAFYjnI1Z7nA/KbQ+bHSwX+Cbx
oTuvguaI+x11rHhc7X792Jkf4iLM8/Y6nN4TpEQyBwP2IMtVmfjsDKr399T0vuyvRsSE4/OWEJos
zi9qzQf9FisU+fyqFa49dCO1qdhru7ihACOo/avEFsvSqE5q5aV6ZqFLsEzvNDIC2ptL8B67qEcg
2a3djdaQF1lCSCVrkHrEEE4GY89KeLYO//7DMr7EW6IdXVzY/RzsrOZ2uuf4xKIcu3qGQ5BF1m6m
cqt1Vh2DzRbyXRWBL5ad6dct4DX18+FjY2dHAvbHAi+wg4abOUP5m1+w750Ow124/yrQ0ifhhE5B
eyRyzasuHl8dFmUKX19m/gYwzo5ntqM4uuRfqS91kbXXpXSBKt4VPsTZQWE156tdQuuBjZcRFktn
7GVsgYPCSskTEXhD0KfUJFsKcOfrXf79R2UngKFAljnefV+jNu+pznO7nuxM2/6lL56jOLJmaTNk
trzJ7uIyhQJbFGXMTWfa8KNPgv6lxCzFy5mjBxUbrWv6qlsVO7NamBjs2yTRnzMqbiBmGy2rIqcs
O+82ry5SIVQ15TaygcGAzbPf0N0OPWhdxiIpMnh/UzdDyXksDwZ/ho84Y5sG32IGoTnxhq85St4h
qvIoPuBVNLOeXvcvXQ+OKvJ4uNiFg6XmFFEzuhzwqn16KWm7xZyoBrgcMb+hyijKCJMaFKtDStDF
k6bkVf/mjH83GpPF5xQ2uy+FfV0UUNhMU/276yg3NXddnI5AC5GgvA+AwdN8h5W9WhfyYu98BMfN
oFdtefwfiaTd5OQ5FjH0qm4Titwv82MEVIFyfCgKOm9frbdWilPhp7VSp2Y6lc4xHn/QcXKhfSOB
yd8JHlR0oLJhTZKuCVK55jffuLbzy7sokHDPunhpz2Bn9s0PyJZ7yoLhYwzEYCq+mRN65UcNsXIf
T9G3Al8PLQEYjX1FS+TrlKR/MWmZYIf3O4B4YHPRbsIWspqmxJoisYZ6Z8kSMjnUJBGflwVjthHe
1ZtsT0YcIR9VdMu6sYTbw2im4pApt6FLyFVl3S7QwV3oTdl4r2cTU1f8cNq5bwTq14VKg0rSXZZH
ztdFHdMFwpJ3je2cOd0JHXLHeiceGXvShZbD3/B0jmMsQgu5MqXKWibeP0vn2xpClaBWs/656NT8
pqID6F3sBgJn9tryvrQT5WYCATcHJT6Y9VGik2GsrPb2Nld+eFn+oumk9m305g6WugQ687XlvLqF
W8y6pyaMw6CwQE1jnWNteI13wtu4LQ7EOTxHORwzS5ewgQoQgG4Fm97OzP6dIA+AXEQXboKucX7T
lZwKfy07BtQ+/c4S7ZHHWfctiLKG/wdohzd+fGqeS+5VKnCs6LMyunZMVQETK8Poss6cDKgf1drj
E1FE0cLrroTR7NUqE2pWIZxtBzvyzjj/44zWsZRtzGs3kAIDhiLcvUCeYIyhcqJzI7esu+gyLmVR
wOyPSJPHCElzBQa/dsiEYVSRj8zc8aFRt9R/0Z5/WS82zZXQdDn/u/kB5lO4H9sK7y/zNsnkel8M
UUj2YMxkovEjUae2RzZvN59LlFWj7FBzHE6OoO9ZcpKlVy4KlI/1ijLxvNHceA/Ng6fOHUTQ9Gd7
W8o9K9YR4FNPjk65kaAOJ5a4yKL+XuOmRbyOp5qqvQ84OmMqdsu0BEEZD0yOR7NLe5GGIlzPJKzu
mDugWsY1hVNe+zmfDXws5h2jNqtDw0X+xrRtEAzgoV/JhgIMXsap34tJCvmuwb9hePGhjo5RazMr
BSlTplvd3eCWzSToa0til6/vv9uZzNC/Vs3MFCHThOZIckRjodIQRILRy6n7Tq/iYt0DB48fVwcm
Q1L5ibd5jBuBMgH1UPTPTZ8+zyp/Ao6hXAScr7p6uOUAsGRphWs9kexOwbnMXpPs4cr7sBw3DjGL
s+TA49rhz3TyVi2+1uV8TfEWmgpVAUkWT46Q+HM9+4VJH5vRyzlXkOT5jwQPQGt/1yxIQPoKOkPt
09pbp94tWo1/c8Y0b6n+tsaPJ81yQzcBZqH847266E6gh7+pmid1u6/TkFhYKqpcN3Fu9p5uPC9V
c5sDGgfJCe1QMS2Vl9msZFHOJpVS3qvmnX2vvvq6NtXFDAtsP9f1FBvzl0Zs1cLsXx9Cc6EuwVkA
Scq81Ad808HYOu+igxhfb5dpsWiS+5QyoMJ8KyM/hlyKrzPaa/iYyt4Zf9rpT1tau0Pgo8q7T1I7
SZsOgGIZqo9G09oWOlVQA94DBE2FM+RI6rXF6VfeT88yC0LQ2SjFVMrlLXmiabFwgrcaZlHfphIE
0o+kkujzwfX7mNhb4P2LPIIeDcjYi+mEwoPqAKrabMIPnIpMkjlEOuMqQfJvWSq9jLm3fUPtvZQw
H4QIgUSlpEfj3s1ADY31zboDNAf6j+eKpYrxcZ86FaPu8TNSCp/c0nZOhM24usD+LoNMRkCqy3+y
mQYHNYXaaXfsqnFVvJPMOj+/OlVwr1UhtfJqKWiahnGKMagCtopkrFyEFtLnGqlI+/YEmQ8lQlTS
EuACVyMn+OLM15RO7EIoFpfTj39dCWB9HCpZlSG/PaL7Owy4CYNsD7/inJIAvRJycOAtqwoblx6e
OuMMsNet1fFF8yGZ1QqnLyPVFY/DATAXKZFX0s0ELjHXtRwQBUzVbpHCLGK9ON2oQZlCb+si9RoQ
ehQJF3nw/grTxfYMclMaZo948MbCpIQh/N1SmyesyLP87N7TEbVPQOY9kuI3yG9YWhAcpPKgz6jB
Gh1/RWW6szxhva8orLLac6sBIA8FItiEQ3gfEIm4SyEzywWlV8pTtgyx4gu+/Tbetrr5iOXykGcd
pPGUSrmCxaUYp6vBYsGYN95cTqsAail7Et14dh8ctyMFyKYAqVA50/EunojYtS2FQ7sTADKkoPg4
/PReGmGWZan3vTo+budiQ0oZkCXt4dnh/g2HzXjnV3RZ589DYV0BLzanMUT2dWw62MUVWynpLsvb
SpoCcJE2kHKqdCmcT7Kdk2UIJ7VwEMdrLJZ6sOKHfFj7dd2H9+339GXHAA46H05durvPmKmhVuIr
5Z4iKkPk+cyCc2iyz8Nr8JT0eI7voC/x5liHiOi5ElQAFTPObefqMegKI1VC3YaPKfXwXnEyFnRy
niPPBRRFVHmu8fcvQZ7aGJRwILUgjScP5Z0NHFOp2rnKQuA9ttSh4HdaxnGNVpLVt3wMv5zeOQ8Y
Zh5W3Zr4+2wILk6Vvtj6BE11BmcTKfkxc14NT0+BYJLrLPD6IM22BBi/aDfPkTNK69zI5D31JZqC
4tdRmGnxshsleoX/8YjkuAKwcrtjzu5LUX5IVoouvN5rPUy93OBMAdzneKCJFIBKunm4bjv7pS1s
g56V6yrWmLnwDRmcyoq/So3ZgWpXxsL3iOXNGGqGruj+kVaxxLl9x9fmdTqMZdUhAjmfSR8uXrHa
EK0Ic6EFHsanuyfVOc/UicqDrXfc8klp6AeyC+OBpKSbcai1TwiIZYXbBM+qoLKBf/QOxVT43pJI
KsDyqW7PuSp4ZW1nqn/8x/68XKrlPUDzYJG2TyW5Ce3O2zwrYWO2h8RzpMzWWw8Sjugh4thutUT0
Ho9Nmv0/NaAbMLUu9P9QmzA+Z5Zj4e9FsZJz4q+HL6LNu3MTfLCi58RXOkr1XxVyxDh4zveyq1IO
v5KwV6CoPdcjewBZEYvPciLYMdgsM2Jm7AEi1tz6N5V2d0hB0lS/191j0StMNpfKjDcqouzj1b6T
5xroXm8ZjYCc0dKJmXHPoEpFDqVn/zURRrohv7tSZ+0iRipfYDeTlyPUwIfLEdrTQucUCUqN76DZ
bcRO44ktJfRQ1wcfeRyA6yvLjUJSUEzEYbr5revPGw8sjSwgLbF1PZq68eeAo4POJ1bJh7lUELjB
gOXOU9Az1V9dHih6xHJaOR2YmwFzoNXjWeA9If+nPVg3z33Y5AwrHkOb8pmMVWP49sbf70O41uZq
KYuKMi8NhUTjjmeWn3ldLttR5kQTqo2wr2o0rxmGH/myujCRYKjoiDnRnjBqb6BT5ofaqoQLJTvM
FSjHHCbIjcwyjAoFdhj+4SVWY8YJBVCPMI5gPlHd/C3RnrDmWWTE6y0VeadrdOAjl2j+YB8XckxQ
7S7NjYzovutG2wxiz1ki5C0nQhJhSZIpu/TeP0KZ+k6LRa3miOXvo92yEEy4KMXZSkzbFU6iTo4d
/0VDdZ+hAw2zdQS3voLO09KsE4bdk27Pa1xZGFV3f2g4gSE4l13THt3WeJSk7Peq8xOFnaaKbnYy
qy70fb8B+bTyPjPCgvmoIIXnASSicB9bxZRjKg5zaGEBY3XXUgaIBPJmt0l0XB1KJ7PLvwzffK6F
RlCt3uGZJOHukhv8DAzvbEtSZWMkHsLlH/V4wu7it2K/rLffDGbC4CFSmEv2HfmxlEsvgS6vCklL
ulPu8cVl06tSgMsw6UVBiCCjxo2nWCbH4JuhhOJVKlX+TFbNorgRRl+i5QyAm27G8ypFbh2NRLkX
8XblfhLTG1cgQJyGAj3zJMFVuPqk9FcxowGpihB74U8H9aUC4BBueUtaQY8/mhd4xSiPbk6M+fpZ
poKZdewilFPCfClAdQTCeDOUOKMj9rx651OvLULImdV+psN1QXtbsTd5FX8dBAyGc3HgZH7ZKT61
DB6oH/3e4K1P86adNUpsjiS0ltCol3I6Bpw09uEGH3PwIHCaneh3MjQYYAT0zIt+cMPkPPQqZRAd
yyP2JBO6VWOITJfiVvULZJUf4yKuELXLcORJzgOFpXw8D2+IaltSyBT4OWWLLNqb4igyJcXW95Qx
LN2BxbwEOF/ragFXT/xYKcoN60uXBMbF3SX9pY32i55vJpTctSNs9tsNrEATfrXc0CX5eQa2OpSQ
p4YXuVdIm6Q149WpYa0QmC5H95ymyWGeRIgSNrsJPJHDiYfWX7jNy6Yw2uyjRA38OCy/fvopwc+T
X798TWhkx+Gh3sT1wFXWtzmynJJrRY6AGvNG4yEcpuk30nq5B29g3cKd32zfroFwwTnn2l0bjFtK
tp4MBxZ9G/3TJCTF4ZOFTYxuXbbZDrRtckL2vxGeVZGMNk9Cz9batI1Rjqb8j6sSMX2bcIluMmt6
xj31iR5X+8VFunGQNIw9GLGBEqOlpl4ww4ONGp70sF+YJ431bk5rnUSM3inSb3+vUyZdNRuneGkn
sUxnSQnz96HS0Ngl85E+F1LKDPDTt+MbuED43wIlYfV2AFkeTk+M0iJjNuseTPDI5Xh3qy8fZGcc
X0FR4YoMkg4gW/nJVjC0HoKRzEtKZmBne76IhADfh3LmqwnWdLfqtZc7L1rOCpMBJWN4p7kXtp1G
Aqc/am0QpLXS37ClUm0EFmATG3IzQFXMNCUIURlZzZdJoMu0Wx5rnUUFcoi0u6USPCS5lasUKhSo
N1XzpuR3cmMd7YFF7EepXwh2xbnVHv3o34b5u6CsJNn786/C0rqmysdb4jewb6MkYRQcJYT9czT3
C6F6cPUuhw3vEXD/ggHrBx8aENwdiXJtn4UjO4JQQkYRwYcHcMVqU+sbylH8ZKbOu8naOSEH4vay
AqvkrPs8yTRbUIfyW4Hy9kIFLmROjIiRWi+hFiFHo5MQkO+0gVJO7pZM6m7HE8t6GjWE9YS0qeg/
fPYK21odo3cSRPccbS7KIMGuNZ+zCM5I18LYQE0DA8/7ZEHG5QwDicmgGO3mO0lL2UodHgHwtooq
ffcoDXvZRJktr2Ou7vkigM68fg7cjNCajBJwtDiRKdadFZjIaAZzZOKv/GnwIklUfVr26YPzXFHe
TW73tbYBX/t/k3tdgr87+pN/esmL+Y9uJC1qMTHu9ChkR1j1uVc3U0zddH3d5jGCfkjG4UbLRovG
bbJyzYtplHGXqjdTq/1guVMwKtLt3AP3qfydUbFCkq3zzdVQ/2N8ddlKV7MB3BDvbfDbgV+2aqxw
2vOG4L8V9rkzmnWiyDTsy3BUf9EqsS++xrYUvod1A7BEfOQ9i8iEOtfXCz+6s8gFoOMAsiWQ3iKI
4eS+Oo5FUHQ83ScsqYF5kocAMFTkNZLSaaewkGBcj5dS66DJ7DPD6JA3IFqjGU7EEt6BWjHG1bPK
TqsZgbdY7fFLAaPXenpUc1N/24EsAcJRX8w0CRRWn4dEEbjXVBFWG9f77yy98NCs5CtXR8Me3Bzz
SEs6PTA1KjDEhqbC6jIOe6HRW+6LaxjkBQ4HY8DtbPGs47QIwX/BetxWCJtW6O1I0rlQu+CskeNj
IxnEk7IH8wVC3tscmMZonKxSFZ4ZxPzgXpxck5Y7iN8bprh0RddxrXSwrfHsiiW7g6S6hVpsyiWn
g5spr4CCUYFEv4QHpWQKKtszCHlICb/p3+GjzE3PG6JzgyYqvD/8O71TFWlmfq8wd3ZxfIm+lvrw
dcwBDdktUlUoymms0WtvgZzbG8G1WCD/aNwc9xPU9L4iIsDtanwQwApS/ypexFHtee1wIr5vZIS0
aDyBRUmvJ31FAxEHUroMJE2MLyBflr73uIsOMtLXgW2pHniCXWTj0eb9vS/xTKP5u1kYPI+Bqhxc
i5kymOENq4sjprewqEpmp7oNyWTiYHQiQoj5Zk4fUdB26DsirqGQTczOwXG6D5rouyyRWv8QP/kO
XiyzQv4Z6NuH4E5FQpT/b+xNMAxS3UgVdYvLFpq+DTXL+Hn1+P6/eubZ5XncLOHa9AXEZx5S0uX8
0UZPhuSi+hXKTxgg7QkhsXMYaFqpC0kxUEOrT8p2MZQrOBn/1IP3EbCeNU21mX+q/xirklTbxW8n
Std3B0dL2VWbGuSaBAZXnakYs7x6qvP03mw7JTIZjWWX+caCt51Nxrp/6psbTYYQw6lHdiXAoBwn
uXj8SSDT9A3MZdj0n9VKtnwtI9QtiK/jOQn2+cv6xIOBehGKcBBJfA4Z4z+yYbgyWfczWo4CaQKl
ERisTu3NB7Mwg3cXy2q/L/35b/R0elJyV5tS7AHZw9iMJ9vD8q6bGbyFHVeu6puOTmb82LhZDZAI
j399+Kq+lEXOiyrQHm5FbQXMmchap9WTKW0ldDBCRCULdWDfjWwA8NuvVgEE3IkrCj8eswnF8x4K
qkY+AH39UQqRebpsSS/byPwkR2qUJiYUzA5e7CTT3jsKGRZg7eBHjpyKTuO26kQFoUe1F7/aYWe6
jZk4YOghpILP0TF5BwhQPueIjdWlIW3bxHJKp4kPhvqBERIcz+gvgbl+rqRmBarWzeRZrmh0EolR
W2BNiyUH83HVmd7YOeZp1mkb8YyD81WXzcfXvHiXPlunVk0KdLEkos3Ffirx4nreVUi8sExfUeLu
ZHSs7a6kvYAwAYumWfPUJI3CId0mnMgrtcIkq5IO/3vC13gm7jCMu4G9GIptcryGo6JbY6H+l2GE
6o7oyjA/PAUxe6ZA6NDR6hcmZgH9/REXm+/5mqedZX4Xqg5+fw+aaT0MuKnOC3AIfcI3iFw+zjDV
ZrCOGMPuUgVDKAwr0ryRhCVPH/GzD0tRbPTgOrZMBsPs7Hf7bG5k02L6uI6f4culuCIIw2lxH0DT
gMjTdctudpXUlWuVWyFuxmF97LCeJob7/j8DpvuzY0zoJi4nTq1nF1VeXX/LcRwE6Uueh3zs6Ins
fd16XQeQYt6OgJXajg4WnACY8f5Mc9KXwQEfXAJ4iZmw9op2fcfq0qX2qE8ySiu629fWN77Ful6G
QIJ2i31iyeK0CIghtRRLwqBnGFF0hpI7BGzprxdz1dKzJ8pVjexF8oQOVdXzU7WwZrgyGvmP2n30
a/92lDA62d1YvGfy772Y4OIimV/SqdXsGe6mgN7A0w8f7jA4btiVYyaXTCLELEzgPhORojKICWcw
zx5u90Xja17YHe1vG/qSBZx0Hx0pn82/83285L1DiBPXqRU69dGaaq0kOreZ4OrUr0g9YaAFrSbe
9RS0BX3uH9sxxXuDzPxXESsVugg1MNkk/iw4QDQjAnW3jr5r9GB4BGitwVtEEUnoJH0NjmBJtoA1
d3Q8C9phTBCGluZE4oFrP1z/+x0DNtMAPkfPWZv7mLN6BRh8bV9YHQvY/yn17cj4yIuKvEqD5Ojl
lbUuLWP0sv19IBLm7siiiqleaxJp3dcWeAh1zxSGsEUxAfCZ8WvUD8y8f0Lb++B7LHFDbGcSweon
7ITcVXa+8x5WirEzQmIFDECQFW3gnIJBLv9REOaA3r6Ofu9BmacZAkbwrV7q1ZoQNih/1fV5Sut6
bezGG1phUUYV6bzEOoRT9t8Af8oz2h0E3g9La+4OxhdJb+werClq+k2iEC+WfMlqv44AjS1FMEsu
Bh+tAUYF3B+VKjoHwmERIP6QxDbOjz9PXys+dZa1mSIJs3cL1hwXjumJlmcIj9G9JGUnpNwiAfCS
0HaiOY4FV5QNKLxdWDvAOlh62+HrsSCnVrovYTHinO7C6r887NWABF0wsCpoh4oH3ZTjkinKQjFD
alif3iJ7iSFUZgZ5wxg+Dk1oZs3qL2u3bc3nT1NSU+Ud0pxfh5ju6BM0nbtEcJhH1VTXeKU/oD9w
XewoNjnwYmLMpKAF/U5OmlMUKZbnKIFGL2b52AqL+0q9PGqwMlIIs5fuSb/P0TM33x1C09SMgLW6
dke720k9XWPBSrgLiSKsSqByfhZzKX6pDz9SwD3dicr8Bff+eAiFEYgNmHxvLGmaZYgtYM9hhO7b
FtTbvJswCt1JiaBQE8rVvJkFFHycITPEwp1jljvWXnOhcs76j0Y3wt9WAZmSYVFiuswEJ7gdAYYJ
FvGaqPubLaQpAD0JGIeDy2nlkHnCXn4QL3YWKyJFP4vauPoCRnlJCE3KEdl45RPisTuEPIKWfBne
YiqGP4NiO55XX+xBZ1taVk/o5KUbJEeLVrH/edSPZD70VTJgtBAFH8/MCGymDLp1IWk1ydJoXrT4
adb7LNgHIKLZK/tPMROYHR5uRK+7G3Lpkba8Re/1FgC5XbD3g68D92jtiw9i9p7JPO9CoJ9XwQuz
RF7RA0VrreXrgpdb6ciDTICx6gGh9MspeqxqpCiKpFXoweqvdcNizK3f21BCTI8Pn8MxsN3jXnFW
jvpZKTH45UaLf59gCG23d0Ou1uIaMI3IPYENKiQBaKekaqRobFNshe6BuZ5wocmnClQTTJQgPusx
259W7vy8zeMuJ8x8tnxeJNowBLOPziteY3Sb9Ahbn+FBVyFZBXZurHbFqYvWhmzjNBT+ndiEpU7u
yywYSDeX0PxSXSaM5OrpkAXMv83IBUkAlHn04wZtb0UN+Unm+VnUSfexiso2VY169xpE7euqmhRO
Hvw80aRZJFo+Z+lBvasjlylO/y1ldTrPntajtZK5tQujlsO2GEZYZ0uUJkd84NRJwnyth17w1a6q
dHlKK1Vi7fn87QrqQMQAchDK0oxW8jy5eL+cSq1sKryy4wtimjFynE/s6uGaT+H/KqTU7d/VVvaJ
SoJIm5u+HGbnNUGOu0zEmVhfZY6CFK09h7KO873ydwKOKqS5Z2qGjdXBaqOuI5dGXxAsgpOdNaMI
t6FbXIo7TU3s8qPVGRLMYxlEpA8Ho7lVV/VjeE8E/jgd+eyorjQlpJXFgOPsUlDeBj1ik0mtl+id
TP1eO+NaSvz+0rS7PI+9/GrnbjfuZzj/BjTuRBf2ReYnIAUPren3ceCYoSMb5YIQemywSYF0rxql
nEc+lO7rj3+kCGvAde9Q2LxhBx1bOJfVSj1wyT+mf4t7A2w8HIUrxTUm+d1vsaVlrYZs+GADn4ha
b1CDBbEqgp/Mfo0dVEoI/tAFDl0lqpvro0uAp4dbPJvhzkx9a92Tfi55zO/2FjMqDAMJEBCpaJKo
F5H2kBmIIUDXdDHKz0iucKpwGwiH1cc1SS8VvGbbsTKncujvh7CNCNHM2EFtVdO5249cuQOw2GOj
mz5DaU8D9gf7nJx620/q7jxZ+PDgDprjDeGVcrrBRFmn4ycqu0MQfTM4B7e5fE/A/B0mH0gZT53T
k7IlgdN99gestCUP/KPXe2MUiPma6GjaU6V/ZjJSO28sWAnR7kvzmTtM1TPVKRx/EXRDbqKAClyz
V3ieLWySREvs14iFI00jqgK7Qz/rPoAN6Pco+NURa1CJkrjglSXgPaEbU3UDgBNDnDfpU0oVrtX1
tuM6eUdMAnztYN3JNpGOcO5ilVpidBYGjtHK7PQzZJ4MplWqRQdBR45x+abBqAiiavxN9Y3Nr65I
RCB3fINPWMX02LZ4/tvcCqVl/VAvReeJQpVHPNH83Dn8EF/+Id/tCm/RlqAbKCeldfWhTETWsXqh
BQvQXAFaKU/Uusk5eiwKd3u8TMv9KD+HHa2xmIaXZpWyOm6rEDify41FwxGxNRvDqq+o3yEcXvOr
3DdGGM+ITL5m2OCbrNKOGLmVvisZ0aZ1RO0qw/sHCs8pUJgFxy0NfiTKVK2RBeqjs9kRWcDlDh1p
IUDSqhqv2E/rOVGfBNGsP/9wcbVWgjeEvFCC7OIlcKFLj78/rLiqeflnmmtJm/2WCLrRAs6J5Gf1
bQJCdGiD4rAJ0I8H902txWYdKf9GcMZE4M8WUH1WV5X05IjyykqsdQCzS/bOo2nB0aeZQFpeBrzD
aLMCbS8iOOi4S+95keod3oeb675D1Arcmq+4F6jCMN3YjvYfNoQyfQbjrsy85DAAkJIPfrPsur7L
xvRDeOi9NeOsc/YC7TcejoywgLMzXilpuFMONO8Mcs2ksVcJH/I+YYaFVVqexn9TovjedPEB4xlN
TtzKBFhA5I40MjZEXxPALbk6Ywjc2eRJsSbz7YGc393AXoI1j/STq85Ca5do53FIoO5BYBbjl3L/
v3iKlrl/WV3eJrgk7ivtT5KE3+Rgs288v54MXUdIEWCrrJQEdrBptrvNtwUiD6UpINUVl8gaMoav
5WPyGF3AESp+MA349edMqZcWtxwan9EJiT28EHBq0430f4hrxzPdk8xE5K/hI/yowjQSvvi5FknP
p4Xz9ZzBT4H0ihPYtxyJnH1wurZjpGaM6ueru9V2YGsUDUK84k4YlBbJA1Ve18r8wFXoAuosgZre
nZSUKTF6HZhAkqTHEkOKgkttc+ALA9T7nIKVjbFljJIpuJ3oFelrJrIYSoIQkmfnuW+jRS5Nhdai
lRdE/7l7r85dDjqOIRquR68vjyvdEVOrwQy9+reMvLxj+i/TqEwb+JsFm707zPpbbPqHsPijL/i5
HBPFMJfli/GVns5QTl3iIWQFXd5REZTszqok8jI5YOFIyPeN9zsBx6KANaQab2nfXbH1I5Ej5yrL
6XZdSXY+CHDoioHH9v7EpdjAMw4UX42CUrqYceQ5PpHkHOa5p5PjxiiIwZgPLVjPn67CPhJSBa3u
9kVYuuacLI2n72Nzox3TrOjwQ/y7/D62n1mQOAZq0KSvl7CdCbO/5Ng7Nam97BKgAzGUTxYdr9aK
eA//XGjV+AQQGvXKuq4U50sCVF2uZMd1P/OavyG31dJlGvJhrD3WFhz9HCDzl/3qWgVZp/J8c3vu
HG1riGC89TA25EAZa5XyGiKBgq4i4b25fKqywuTGhOqUKuRKMg7nx370/tN9PAtcRH65ItVXIs2x
AssfqSPteTt3vFANeGh5tWrUfvc1Wk4IMuFC6DM2dQJlRwEgVHPGIYN78QZbvMk+uY2Yr1bA//yX
7BsvrWCUIFRBZFNN88fs3rHZa2qsjxsMvzhZUQTxQOWj029MBMooE3eX6gbzTGqkWn/f/j/9zes6
a4x/3P/VAQaEaLJrYJUlnc7Gx1c10cwGV9R5fFNsQg8sPaE/NKvsFsvE/OrhBS4jaW29KtKj4rOA
myFpD4MHpFwjwLtrrAbrJBuaoasMjMcDEHxUghiMQC9iElJ9lBCakyZq5vqWoKcNMj7oiLDKlZEF
VrxUaZxCq/UrZHbB5DfSlCBHbJ/noUnD0VFPBC/KdSc1mF+2t0RxW1RiI+JePQEQRQq5jfga2q3k
/OZjGXBVs25uqE3RY7nqs1ccD6tWyl+mMa5p+MNPz7vie07qc54xvMzxI0zdJC7qM2MVTdoX6Jfu
E7vWThPJuFmHAnE8NflmmOxgryU86nBUfpqx/4J8q90OtqFu6/Id03GOpYgwHV/WmmBH2cgPaLHn
MbAjpMFhDgu8EOhVOYBn4BHg6UjKpscIcu30uVmalDFiBtyaqMUaASHX/mhwlCxvpGAeCGy4pzU0
M4f6bAHd0N79+Wb5RenMYiYzbyYyefakviqgrZYZo11wKxF6DJbKgQuSQROecgjqX66d359WFG0o
/aNTjEVF2yap8g+FVSi2FWwCiWrzdlOdScJ1TiX+ttpO4TI2dzdLE+exgiEkUiOQYfUbqS/yPfai
3LCupIWkZASTDo1Hjv5hgt6CSn4K6lRXrglenfX4RhM+2CGvppqNYTms9WnQiTF3UanTgapPs+Il
MkiO6n3Z4wD667ZWndt5Q6e1HlEohTT43+2Z2R9HU+bjpeMuwrG/zd1Cenz0Ts/oRFOhNAezKfPo
ViHYjdu07Imk4aqvJyNRipVEiiCfFmJlXCtxKc/dlr5hUyb7YkfW88t5Wl8dRp8BG2oRjixsu9VF
Idgu6z+BsCsFX3gfhyuUIyPb62Qfnfk7IU2zMnKS+/sx5aLoUg8pZqVkyLZuq5pfR4Xm73SQmC+x
RWeZ478LXxRhUdbjRp5LX+Kk8wiBZoNoBMHLp5cMDQmgR5TBdqAY9G0w0Ie+73Coj0rKx4KytNmt
fh5GzpUJZrMcp4VnsiMTac91rKlQGNeCOJzGHc8M5tZAtA4+miKal08f+o43DWS60VB5XoTBMzEp
ViKSMHSBVbXJYeWizcL12NKjyfJoqwY2XQrL5/P+6zx7K7F9kCWRePo0tPBQPBmi/VmgpDjyxRs1
4WeK38+n+wycZ8tOTHGZN/aIoncwupgSx+fTSoIJ4GzHVGDGg0o06tQAmoOgoJox1O8mLXI38ojy
odAbToQlg/fz+fZ5XKHp3r687/dudqqKYfr5yIKBpAr1D4+PAD9yfBly5oMrgxS5jfVtn1G3zZ/U
7G4qGxF+ekw6uilAalktvMBpuUPja7zctOsgiU+nrnEl3m8xJifTOXT53YddWUsf68opzLSEoLWp
fEkb1G0IEG7xC+jUguVPjK7b8j1h1iA21Wj34il7zhxOxWEqlSK7J8RAfh0id/fqLxg1N7e11881
7DFBG2W6J/9zV6h/Xyf9u7s/ezir0+xEHkhIbPIeYetGdW6ivK07QUhgE+W9m7H1YnmkFKkwwbYA
dF47JQVElpEBJHek2AS3K2cHacBKl9FZfs+bt9sTVgjO3+42ZVQ5sQk3Snmpz1U0dpzbD2d1vw4B
iPCSSV7iSmAuUpw5bqQ7+TYoNEgUTIKH/ZolLdPAGl+Qy7yvEjhm3zKo9XruBIWDtqZdIHo1KrrX
kjwZenHWXuJe2Ylqb4ycAgVYYJpu0EKfpFEY66lt5OlVBTZEFycNV0FRi3iBIWVMPkX5BzR+ZXHC
Y76K+CxKnxTWOViqfADI3T9fACfDUB4rgOY/j6qy1XFI5y2z5PJ9NWVraDvGo6TmCRlEKRIelsTD
JIZu71fzBR+m4k/VXD6DcPpqIu4228xXyeKRCMLs0vziJk58USfRMelA6lmGwbuUykakC/X/z33y
LFViUClskz0iWE9SycAZBOxCHgB7yooW9bhRXQqxEFNDZcfPdzzZKESBYktlKX2MAVm67D4I61uG
g9RBKgtcMtTon8lYkMC+DGWeZ5sCJCdKBrJY0kvruvRQHYpq+odBVZ4RaoGSWRciOaPxbdF7KyGi
OOCybYE74iJReP1ON6MjpBz8ldGkyXaN5CziXYA5jbGJg/U18SeiqQSa54NB6bZJy6LZZ8y9MqwQ
SL68leC2LdoS46sf02QX8p7GBt7s97I8DOf7Iviv2vZIW7Sm8YTvELyd+gaxjGVWQPl9luof2XUy
+7pLPAU75Yug7v6OvDdQC+6ITtvf1JeaupYBXQUjZ0oosLSbJtkf1l5iTaz7YhjF90ozR6ejj4xF
kL88uJ4ER5VHp61ReZI50KMjZTds887DfDkI7XJGjIXPOv99t8fSo82oCi3BgxP7nABLkuM4Gc8k
nHTTNOHXj/oFsogaaadcW5a0saQ61ZDvDfCLoSluXbiGwJQmfI2g8dpKOA6S3mnaFKfAgn3au363
5YPoaf8EMMN/2HPhWBWRjEZ1V6x4CQbF6zp7W7V3q/yEXtWrCW8Kk3JGMIY50Q1CRVtg5swXBCLz
Z7j14iWOLlY5W85HWy4pu3WSI2ktXGB8FltKGZwqv9Vc0Q+dvPPUKACuUohfwsSQkecmN2QisAjZ
7/G5KKUOeEO2KTeZJhhxnA4abovgqjmsCnT24MKlnOEmmNR6IMJhF+mNpOWO0crj23cghFjwcbrS
q/KdFJXQIFu0NGonJGZElSF7EL9w3y+SFJkPRleX9HZz40+XBfzYfmwogJWQ7u1PCflDWy/zHFWZ
4l4Uy/beuMYfXtqkl0hPIMlmyHQ84mRHpAik+Qa5va7ZM2lsW8lVEqiIrAWADzcTreR1dVnECIML
eItQjrg536pSOE8gAjy/FaNxEzhMhgxWeR6eoEkzJ5C7X7qOrsBZFcn4sBHoNrCZeTSrfcKURT+P
yn1Ggz+amDuhNSz+sDDe77DaKlbviXk09iL4SWmSSiVfIg12T4JhViDCFG0L7pXsnoHXiLbaXtsV
yjVjC2eDTGqwUp3kLwRvCmc4DMd87BjTWQJIyVQZHljIN8/xcL4G7rNom1GOctI+YaBMZfLBqu/8
SPmGXCXOfSEYTGRhzFTk+E+i885tvegxtqbpnZq1qsyx3rP5PIhQ2K1UpYUkUwenXH7c8W0+JyTv
Fg+d6CHIOGvvYGbfFNiup0lB9hHWd/2O4yN9zphcA2lNNtEnrVFJUYYXw82IomPBNPXTt+//S5nw
GIt8+b6Od3wR3TlMZKlkyF5eKzB6+JHpG2Ia3866Yzudcx0Alz7hsRsRKUmKcQ/4QlxI6n+5zSY4
/+u0aWzs1rqp5/X3+Y1JZYL7AP4P8MFg3FXZoWsZKW2nX4LuEMifCwHXVxXDiry64sucknD0BvVz
ETnaTg8OckApMS9j5kEyDrBimhFxW49CvxO4z8ZcJq56wRZbghOagaK8DkVC/jpGk3qayekS/V2Z
Nix6rlNBKghDsgKE+65IpaUX7ephh8KpBQsYbl38dljMLc7ZoOSKr5kfsfDwv99dlu4ctjFIYLFo
aZDNaxeCHSwlRtDCFg0vkaTA4r4ZYMtHW34ZVE4oYsRlm0tikSkYuPcKWCPxLh0Eicwgm1SF8uaQ
65lOKo2WV9jfWxc8QWORS4mr/UeuRhxIIoiDfFg7yvW8rgxpM8u6qhQmJxOvJkWQ1Y60OCaxlXDW
k1A0T0qfNWNCQYByjpvmG3jc0nTb5fY5qEBtj8Tx26mtBnuUarc3kuk5wLU4kcDUmZDBpsVBijer
PzripScJUhhcEmT8Petzix+fB68uR8cTZpDBghD1TXrtg9NgkpbwaV/+Bo2hrdy07MbkhJx9gCqJ
+OEVxC0nzpKaVWLl3DXBRVV1xGTt+/7sGg1Edj0kiHpBrtow6dSmLvdi1R47YwUNWagyqsraAuda
wKYlFx/BNJrIOT5w7hmlAToSZw35DjeoPRYY47SpZkoPGlCMXMRwR11jKce3pspYGiRbGQMGMIK+
y0WjgCosYEwIomnvsKIqKCmxBiD8jn/7P9hbCYvre9Lo6lp5LeD5JqD0mQRo/LAwvXsXN1zS0gqF
zbU12wJhQEEOBz+PmHhkD9fT7LZWO2D8hLcgIpoludJffjXzU2w//qx3TxeWxsTae8g4xZ8QV5V+
Uu6B1Z922fLGAqAlMxbZDcKRR0GMyZv0DsY/3RF8qSEVF266EmlX6hD6MYL/WJ+HERS03G8SBOhu
lrvUZ1gVFVhL3OpRaTVRHjZxxN/Sr1wsEpWN2hmhoWPM97ln0vaADtSCg6Xwx6BZ9ZbmDb0Mlzw2
8LS7SqwzjaOYghf36imw1OEkJkMOyhKkxKYuFwF+t+WyUlQZwlBgSikqZBltF90ERtGcOq63NFwO
qJLXy3Vug7chPWpryc7Ap//b8GJP+YJl/+T9z9z+f62o2D3lB7WSMCw6U2i2CMvXuTOc5F3bb6+G
YzInryUOr3gF8OmQSkl/rdk/5RgeUCs5bwrVXlpFUzwOuLpHXuaw6EhV2Dlu6tRuPBLuVOQt6H0T
xZK/j2m4JHxWzYrN6K1YzhI3Fz9Fi9rJI+C7ffByaHP9TeyBSmLCqauUH2MCWR4O27jrdQJG3ECd
kSCrSpNjn7ymgf4yPMLTWBdlGm+H+p/iFGg5RQB+VdNn42cNZPn14NHP0quUuXKpnR662Aus8uvi
qA1DNb/nzE7P2BcztZdoEpOtlttvOn0RFHwJKyZPFWxetAuNIuiUNFNDYKi8dW0bEpwoDGDZHX9Q
/e6w19lr4XL1ZyTZgPNbnc7F3geIlJlzbVinQMbaz9wY/ffZ8/Q5SIvgavQtTWD3yRpizydw0x5C
7rV5FUDB5NUkUzif1uq+XBb6PpSZfs9Vd0xbhzL2ecGQtPbfGRebRm2WnLyctIITFagzoCCcdKLT
x095uMLLsFN76C88+WwRVuSv1eiHJulyNVewn8k2w09+V1Tl41ro8YKZnp1YUp1WZA0Vk7OmwG0n
NeIjJ8a7RG4F3lVDPB9Z8PQK7/pqszBq4xlUj3lo9Wc1iJShDMwNsFuoEobFIt3spQ2XKJwZyjp2
7RTx6gkFf5+BIKAOwEsgH0TjoNAFurO+C8g+19i5kiDrMae8vd1+ho2Gh1ndSzoVhGqB4FWjjm8H
QFa0Cmed5/S1IYgbLPn50XHiI7Rsr85MTp3deqHVYWOok5wkiBAnY0M2MyAeSpMSEJOIA+tJgRoL
qqhUO/kRGGYld7nrkVsIrjIMCY3rB9KyBuKvfK5YcEi95X/G2qc92nwJRReh+D7qEc1HNakkFbz+
q6B0p9nWcu3gyadx2LltpV1ZQG1bWYr5JImXJvi6chGHw8s2wX0D5bahean8tLL58DfiPcDDDho9
UR0SnFR9/aJsbqK009PYrjq3qVe0H6hWJSsibHmKq/ypbWoCf9DtFaghQogagaoV5yIn8mydQFsK
VnPe1cMJvSDspJGGFf/AcCCXNNWek6RWoVe+zNRJhuHbCkjugetTI/OuBWu0YFn9AKHXClIlINb6
KFbHeF7U++mxPmEoSdw9Q2CmuYTwZpHz4iRh/s/NTM5px3Xgqhp+m1NnIjqhEOc1Clh6TKEpKsfA
37beZpsaWzsaI9SskBaHkZFOMJHZRNatNVU8pLk2UeVIi2USBXAaU+EtatO9OZyIkxvnmJsRanCT
wxsxKjeDxtOJtTQO1NTS3kuGLXqYQSBJT7hiYuC+iOZWWFq4uQclpHQqA6tgTsNGKm5n9jro9GXk
+S5f+lc2gPmHjI9+IyzvBDN10AAH0tpRcdRe54JUe7czLdVLlZ1b815j0u62BG4x7/P95i39MdLc
UIcZWF5DC/XpICXFOM12SoiMfSIUbrJLeXsFPQPkCguSXjpplSghAS2Cp21l/S6UgPcR+xc3TxQX
d+cfA5mVbQUSW73bmeP1Mj6wb3HsOgidAj626Fzw9WQn7EwhR7tlmZob9cBg5y50e0yyEDu/WRl9
FsziO9ZEup7fVlrmWywUccWbgj9gr124AnGCV8B5dVdLgVzEcVPP0MfarrEcj3TAa4Lb3z0IN+92
SXZjLrUg5znBTAgBi5xe/Imb7RQVOd5Ks3/Ou90fewLoA2GrnuXkPXjdv9PhwYOkU6wYoHJQ3Lvd
fMeIIFTVhiJL6syIuY3rJwvxqk/h21HZXW828FCpblszRf3wId0iffkz8xGLcAeX9ldTLXsliuCC
NU3GrIdeCoYG8mXRMbY5AE3n45PoMIxHBe4yL4kROK9IMByRZYzec93wDxXyLgXgGPbzZFShw7FY
j+YUEkUzA43wYM0V7QfIPRwQbyuws1bCHodA9P885hooeaM/4vByhin7kftvxlJOb/5HRapRg3V3
wC9XVw1EwKwHvL/OpdmqpsoE+lYyMu0Gd29Rm2TeOENPI+Iaei2+kHoKTrXUe3NnlquGCOdzXDsW
4vSa2P7q9JMHFIk2mBP63j4xgcg+HNI4gdkhx/SAR4NcrmxXBoNyOUZJznEUO61oEAEZNBMJBJ5m
N2WZ6Orh6vok9QG6l7FB6qGp0ohWSjeXikOaMDu7UjeHprSen/FgE6qywZxzZ04g6xW59Ea4S3fP
qC5g4B3jEhQG1irZUVmKfYA3YATtnzgw0jPw23xdzzP88oh8BOqLjE8HEZ0NmvYXcmf0C/EPU9iQ
6P9XbV57ELOarwYtuB42wujPmrK953P474Ci20emE2OdL0Nea5hSZWxGJ8mtxuxfxA5UAIEhrTfO
FToaFRSGUVff/9FocH/4BzFz19CcT+cEg9r1fl2EtrhIO3mbVUtgW3Mz7CSstRvE0eRlU0hhMvgU
5S9BVfbRO+CsKxHJ27cg9EMMSHEvoU22/iPcztvUDLhN25PaqSP3Rbwwl6VXJA5pzUlqM9iRcZxf
ksagP5/BYGiIEBtnDEcS47Zvbn5sgCIjDzGsbjFlnbNs/ClDrrbIwYxDmV26t4qTCjtbhhxrDzOB
fafboPq5DfYaESY8ySggMHAC+yNgg6T7exu/dZ1mwQJmjy+mWQqtpuAe55D+62RKub1g22jYBkJO
o4It4Q4/67J7PBzb00rHr60VAJPk1Lp2zbxN7Rw817HI4GrkOGN2cmmx+Znj+8KLikYPrXw0z3Rm
dg+eiv16/5ZOzgRSFVW6S+TO5a1E458EdMrTIXlgwwJ7bJa2uEgUYPnrl/vvRcJ+bzwmsnpbjEq5
0F9QCa0xx4UUtEGfDiywHpQktEGQMYz7zLNAdYlpT8AllVhLI5XtojfBmHHh0rVyXWXD8D9EbgJM
IRJqvLWNcn8nqZBLxlxm9DfDSEtY5ymxK0bG/EbK7CKY3mgqhF8UQzSDUoScwmsYSeQE0rB6kFdT
RP8Z6MXBgPtD3jtcMHD+2O8frZf41STaBFPr19dr29MfBBS56mF/IRUfb6y3F0rVb8UyjUhuhPsu
6nIV75/Xta+61OF5YID7N2uwCV+XyrvfPjG6AgNT+MyEWSagFNcT35CnWkqVGS3kXARN3I5GJYkl
/4zBt2tLVdZQzqMHxlRL52pZBY/UaqUe6+C0YNGQt/aFI5Kd05RmMv6OvhTce1sphsVWya0Jlo8d
rMRTqgBDnHTaS+gldh7negNHKZO0TP4AEh+8wRwpNadFTh5Aqx+ZjuEXjdHKTI35SVYvaIHMB6K6
isaCa3WJV+Dm5aL+FdjFZ40pQuvuziSAj2FcTgHc2cY+g5APvgYwh8viLWfB5jGtgr0YaTJI2MWG
Ts+hjAhj9c1LaLo+7vIFyv/tkmAWmjOr2DUOCJPdbF8E2GF/eNAHsOWJ+ZYbmWxOXVB2iz+UmK0J
Ooex4iatnJzFEOOxtyX12VPRMJhkyhUACM//XHRQDSijnL9snW+2EgMrd0q3UDN4ga+ANRzE7mjE
lPBoiBVyT3LZPYR9mPgYmGAGaTZquy7trMjPqbgOzzqmlT5SF5oVAAYp3qbKzebpOlb1h9ZnAXLO
TSiziZ9FXfTZYy/x4NFbNLBfa4hJJpVN7JoAEUn2+dIzBDOwa5010e0tkfIBLydEkke2YEC6l4Lx
6clYbuYNPazXQlRVIzJB/3B5jENaVht2dY2iE2Vm4WEFJoQ52EyebD+l1XDSb0equp9k8ylSnaj5
MxpoVwQZsulEXpg1PhOO9ll+a4y1+SRBAGBMNw/j0brbbm6x+cepyXjmE6z+wIk+vPLQWc32quoF
9D8JRLOrzKOmthxb5/vaxC0iQWTls3RaxE+adaa6gL//kGANMlWflOVZxh/V1D/ZDNQbpEbHH1Wm
o0ws7KNzUJji+tdih9fPAdsjYmiWV3al0qFWmJ+FE/wjRaEXWlCKyQhIj4IdwL9/TkbVfk2EE6Ck
nFkrbVPSuP2HCsJe0rHkKgMjYF/MVcF1WeBugjjpCu7xrlNQTZ7pwEDxybTcy+kfYJTHay9N3vTt
MDR05rWJR5Zbf3qjO0MnNr2YSQUQe/srb5OpgwCjF4yFsrCujAfZRw0sK41YIk3+DFlssiMjZYHS
GoNd/mQ3t/pR2rqOmh5UehC+6qTsYh7tHVcYYLXpwSveIMDfqhoO076Ps1XJVcYZkZg+kTUT7MQr
+wtxYCgwmZXEeUxU+jmM6bY8+HlXJ0P4eX7tP9sQ3F702FqvKGXFdiZUUo6yBVKDhG3TZa9jQdLz
AD7I3hK7TDJtxQFloUTKfDohzMCg4czCS0Kd2UB1QViMqSTaX8mzp1xDfwzY9NnSJ0xZOpCt+O5H
ULtH9wULurBU3jMOMkSI/Gb1QSqR/DMfi+cve62dfR6AcqyKdtCsof17oCSL9cHPX+Hz79+ler8z
nKUrKKR+N18fcv3/ZNeMOcoVFRQ7FJrQnJ0Y2u5dzDpcsrZJqMTgk/BxLGMcyIPm704tjz15yd5m
AnzNkqGL3mEj6wk2nf18jyIYm4KrkkEgzJuRuyXcnlTUoqX8o9OOiQ9zJYnC6Tw7SHgtL36J9XmW
yuTuSU2ar184Is6D1Fyyn7veNNTNypHMaTZUgDi25eX92bMSlii3kkxSBNwDPMl0VajVa/FEDNLj
ui1llAVMSZchTA//iDFBvriK7j+olKa4OPbcfqA/Mbg4+izeKNLyGIqsT2gt7yyqcx+wwtnavUTD
Tmisz9LC4QzuddIruESTAUFgdt+mgIModxerpp5PnF2ID4yjCjc72mCRx/lS9ghdn2NuPiZLbu6C
WWCTNkpDSkwZziIiJDpHE/WsLt1Km+tZKWRLFF7X10kIe0+Sy7MdzMQwPBM4VGf7GN33eYdIxB72
NuQ+JxnyeCRaCbvs7vgXHyNe4c9gg6mbeAlxjiitK/5VmLIpPRpTfHzqCjiyz+nWZvomvOHnlCew
05qJ0jIsfF+5it0LA888W6s1+wg7JycpKfgvrJC0vm8Pm2Xt8vH+oRbvCVTGUzTvS9wjVA5oB3XD
2+vtPH+wXM5vYwtztFLfDkhMINm8HaRojVq8r19p8XzQGxp5ysqevRiyyXN0dkJetZnaeYDG8bsJ
QyEFZcBtZckYOzxTsrVP1Li7h8n/9/+JrLKVM1PFb5DXS+lVJaZzpgiAmjkSLaZsYf+nCKxueqvK
a5XXZBiUZtNVU5AwnO/AypAAmz/Xxah+aj1Whmke9xE3X7BH2JPf/gEiTy6ZLnYz4ttu1z7JE/Lb
qm5pede8SvDmq8nJekc+7WyxBVUM6tcXXb3mq/5PQqPO2R96bR0ZKbWKvEqYQFrVJ7kJx5vkO79b
zlyIene5M+hCIclwK5/IvJ8BfYMx1armgliEjxXUwqaGDESBF/gez73maz7hce5Kly/3Z2oc/OBo
O3OKbYe5CLamOUMdWd4kxnMT5qWHPyfYeZsjpsDbmAG8s0vBgMrZDau28TRr2yR3FSvn/L/FceZ3
SDGqHHtnviq6MlNibqdE4Yw23ZLQa8EepS3afpjMDhx6lt/8CQpVJ8ylH9hvGw5j7gTn2N1B8nzx
od0KlBKvlbdPwJm6vQkEyJRBR6XvIFHdLUK8y310hPc9x6vemCISq+y2E+GugzNnUaFdvwLZJ6Ku
YBioJ+pBzO1eCaIKAnbMWd+beTU4yk1cuW2bFr4lONW9QvfGSkl0Sv1sqlByW8KKXzwr5CTfjNZs
+ZAuccHZ7SP2DxFnupS89f7j4Dl1wRSieV1qcwPI77PUxhydDDwQ7Uw+Yo93Mik9z3Y+38A4M/nC
yB0GMVhzksX/G6dIAK+7jNwcmbbxxARqM0fD9/JSlYp66hdJcrg8LMoiUz+sEvaATbRSI+c2twZd
OyoVrOkPZVZ5q67GTe0HoddMn9aiVDRWOPTi8Fi0vpmvND1jZdsk3VI+QYvQweeT6WQKXNS45N4X
QBiHWfZbbGBrXgs0m+jwZFl4kPj5VqEskzcMBIrFVMTjEnyPiobQFPGljyTwS6BYw1LI+CX4P6ku
BEjntl2sd9qMdLUbYAtUk13tpNHiPTppGSVOlRbPNZ92e+9o8vihNSrU6Ysqr5X2V1PJ5X/aG95k
JFWcG3ShNqRFAKMJDBWrh16pfqtHx2oimviPuCRTBNaQMWXouFSVlpr/Nyfh826r76Zk8WOk/qET
sXpZRep0z9aCuRGboEBnBlocYX62mdWup+D1Qqq+Zm5ahMhLnXLdib7xq+2H0EPUjjFEZ+XVRNLV
E4S6VX9fnBc0e0RLTQTyQvHL2TClItWpz157zJxa8A83IdXsV1oaD7sucIa8HwdbdZt1PEIDPAo0
FSVc/kXnDcf8l06PguM6b4VGygOXVIs0aKImr32CRnIB1SWsYt6FUl+Ce6nG+ncjbniatlvf20SA
VK2x1NKbfYXAtn/f3x3KCDS9MAwSspH60KNRraIFnCpQyRyIiyN31UxAQov+V1OfqRGVDMMWHsEG
g7fFSpY1Lunswn0QdddipKnOjANDJUj/au+TbcriNaoiQ525FrtyZAoz7lHIT/59R6zSAh4uvvxB
UwmBWRDGgFFuVYGUSWaKu6cu6SQJ8eY+0svtigeiPwreTZn1aOVv6GL5R3oz7vtlDkhsI2WFaohR
c2HPbY/KWkOtFwlB6tgsrYpxRPzBlX9Zfeagj/27ZP1BaUIXHMs2QwPu8AoUarO7YZc/WuXFOoP7
7dSPS3GGkHF5tUMHH+MbiJmRtTOF0+4Q3DHpO8Hh6P4Le41Q9mlQRg+2G0diK8TAe8aKc01zDTTD
uhTAlB/HffQUByhYM2IBWJXchHrujjFbcvOTvse+nfTaeXv7Z4YtRrIMpOUgEYzwJ5OKyiHA/4WQ
RN51J58Pp0wMiY/BsbDwPpks8AzuxaALu9n/MCevIWEUHYDMoXaiCoYA6f4KZYiIUFETIaUB78lz
o+YmcaFAly2e3Hd87zAq0vdJuP2EaG5jopyD/C/AFp70OOOrrKKiRGF6Oan4AQqlJEayEcHsA4RI
3pqIo8kcKVb2D5fEExsXdLc+NqBEpn0Nf0vWvSuYOAAW16R18YD5UePsRd6gDujKvtxhLOaUZPBw
LbEr03N9R4Yz+bSy+YgDSA4QtBTvYd1sEbIvhOahVhCx682T1okHAIHNtzHmxFG6dSDz49sXTTt4
cSgmO01giD8QDN5cXcqoGOkujNuvGQtXQfo9KsQ+avppdS6maPVYpkZPgAzev7E+LA2q4G/c4PDM
oX2AdjvEY6+WmADEXYOUjsq59aAB1Z7VcynMiAu5LQsC4Pn5YlWUii2mo7HgGI/A9hLR7Rde9RNX
irnocVDIkC6gnCLW5vnTsQ0rM3jOCxCOhYCJWXckfkDQTir8dYMdCEaKQyzOBSMar3rM3JzmvxB3
Rpp1P299qN79Ht5I6mVIB/eCBuubGqyf5Coa+tkI8q0vxg7TFQJbFFSEpJikHOtMUIzJdp6x1E/b
uzx3z82A+yQW/3BRhX/BMsp4iyzIggd88Apwxftgx9EIkhqaQrXvlHIpon4UhqDDGGRJDZGQDA5/
Ku8mVnGaT5eIrViTItk0dhUxzDVdBDMmgusLW0dyqeR5pJ3qvpN4UribvrJsBGBbDQPlF5wMZWdG
fjVv/6UY6bfQMOdgcWL3BCbOXqP3/lhkkOSrl0F9KE4yZSSHX+9crgOAFq2FdbF3YU4rdfHxrFGH
sYFebn96ROoPm0gXczfLc6e2DR25JZ++T+yzSQ4ONcZFplCU3zETfuux4S1cAG8rxET5OOD5BC1i
JSUwur1skEw+va2GOVd3dBYaiUQ0fTFoVHqDtGGKQq+43t/oIOyYIv+Ga1fddWS2GJ5JuY1k8KPH
iUSyBjpNuaBv7oeS2lQKTr3d+Kg5TnNrxooJhhEfYvdxsVeIfmLoknfdtGbi4qa89lSdHxivoBws
vBMvF8F8bQmN59WKlT4hB6uHB5BzjhruG9mEH5ld2i2c/45NdfMp2s9sAUieVl0auMFld/GuPMGt
rNwuel3Gdll4XMCNbWG8hzyqSFF7Nd9jATWN6I6v06rFc80y0Sn/DdnqiUFbfIz3yPyTa7Ko96q8
p1GMGe74yJKXr38eFZLLcjX1AE5to0N+vbwOy9zU6aWw3c4HB/dxijJTuRezJpjX3+f6vzi4BjRI
ybv76Iud/asJU6megph2BI6rj3UujylacJ1OabxZRg2hYaF/DVHmF6E3Cslz4V8wZghR99cKKru3
BK0rXDMA/fBle9EH6YqpqsVN6NIFn4Hz0BM+/XmuowmnQ21T94BzQ8uU9Rv4MK6NSdU4OoAINbZJ
HOZlqQGe9vqzPWsd1QjZGJm6Zr9JPSPzf0O/ulcTu6Hk62UaXOINvn9O41k6hkJt9moFllqcsInC
zZFIEh/dWnF82F3+B7FIwFWjxAV4ppuJXgpslh6JKM+gljv7cHuolCuvxTRuB762KaCIVXtVB3n2
ovUR950WzqDrqEtlo9BB5BioRqcEg05FWNUcDhmUXYcctGVNh7l7yJ1fc2mjmAXM14kz/IKzEOnF
q2SkiL52me2I4V560cvOIib8MAe+ugFieNsPYYfwY642Q0Xoc+EUz+/qvteOGtUfTRdSUoyj9LgW
KFmrE004Ba99wI9sPpx8NVCP8bkQ3X4MJ+Af9HOOC6Cti9eRRLEhQjGhIuQJCI9/1QQJedRWAA5U
FMXkyM+3sSQzLs90c7fMCgNjNOaa5OzNnv4ZVCQfe6ikM8anBIeq+qcgUycL8ejpfHnNJr4NKuH1
+QuY8aTN8oXlayaxNf+O0q46mFjXtinT8qbNmJT8wtMjugDxmNPzteTXzM3Hqxi0d/n1wkrhwzns
Ue2fy7UA2Q2MUdnPORtH3SqX/M4Xae2Vd4SiaOlQTu3yBBHOz6npvUisZbOnxtIF7srJoDB/IVyj
4Gj2Li8KWWEQzXWC7Vu36rG0u2Tc/OupMmXghQgP/BWCZt32FeFGKvdkmD5rDo2fnFVBfUMBpTs0
KYqkrvUchq4D22zAV1J5nvum50NRRPA3Cyx2vT1ffX4o+pT5mblqMTvSLwB8sY+IYpvVUHfdBuGd
M96p0fUmTSmuCJlMAKcTBjF5xU/9RqcNJOCV9FgAeJ+v2LXu4lGuMyVSRS/I4m37qpmawAj2XCvr
KqqfWtk2r5Uq1150ocOncQ52oFOd6x5FFhtj7REc1zdSjCcn1/Uye/q+pC42m3iniFCU0vfDuT5n
GlxHqyctBfk90YmJpG1CMUbYAF0rI+5NULch21OFbosEdkV7A7yJyv9NAiYTiZ5f3LSiZ4+ZL4hv
yIaIjn1urY9dcS0jlAjiaAv63zf7Ih8VtXvo5mS6kXrFEJtWCvlG+sE/zW5zm8lZw9HEOWmMwgFX
MSWYDJ6k1mwXNh8BybElKL4TEYkwDwHO0fuzY+4ALbWInN5GD2SOwg318Wb0QwoQR2KOZP4e1cj0
/A1jWloIHVDbGYxGDdUiuZBxU3EFeAv9UpHzjnjCrEsciI5SG0nwp3SUHJhdsh5CQcHjBuZoROaX
oFlVe8ClEAas7SSyV5JES6gOMBUGfivExgh7KtT4OyIZfV/P4ViTWq8kqdpOK5fNWnmQ7kejysKh
LeXdooSBqAsyKcBkraVoqwtpG+L5yoG1RHdNdg3fWh4wS4KBScwAxDvySQsuqMA9qvgBHFHjE9bA
W/5KD/a5ey07LIQm83P8vWK0WnT3xUmoOPbEwsBMNuv7VH0QvWKlIFRigkR4gx+4mzjGwB+aheWF
t1YFruuSqaxe3cHEdqQO6VFPDDOFH7RBKm96PmW1eT9vz+Yqais9HyYQjUDOrCDaCoFEBO0fu8UQ
nHLmqLNvGY/VeMckgCZoCB4fPZWyj4pGy0los9hSJKegKsukdnGEr/Ic5rA22wdhCihiQgjceirt
Smja9YdWav5L2vDEPEURYhBp2DKG2xjF8IcdaDxZdIxziYxFeQneFGt40ld7wbieTSKUyzb1Cp+7
diiEU3uj4sS8Ipl6eHL7eUjvzaAvKsfHPu8MD/eNGNfV66reDaf5IryMXHqJABg9hH4wbYuo2MzK
KiSBItSgdTX1f1P1E2J9ApJ8iKSwEBJMIB7m3W70x5vFZbH+QVu+H/G0OQrYlZPUfd0sVxTQmu3f
+xLm4qxYogAprlOPG+hg90aK2+hYfkc52AVdt5wOD7OXZd1+X7qzDGsmnkr5CqEs292EgaoQ4j53
MxUWcHsnqQHb64wISxjkAxPei0R9i0njW3Q0mdfXD5L5Alhhar3wOgDU/Kn0qvenMkglIQFfrMUD
SR9obx+ShAr6T4KloKITfybq3B4z2OFyiiYYh5NyLoodPUGeoSEjJKz0BNXKRIQvovllaPcGP1Ar
cSj6YQZ8/K7KO2wfvT8rj8AAzTansLn+TeCMrbcGS2aITaXHFYyMqTKgwCxTNdp6RU+gCekVIIRj
0YxC6NyH9i9eRVb5PpP9nnW8W2vKkbkZV8jsTdgK5qBI4xDuyWYy927KAPXu2H6s6U2OVTHPvZQ6
edAJcEq2gjA8YdT0GoCel132hI8jmETbnBErK0hepsvjZGf0heeoonaaU5Nn74RcI+UZU+itzvMG
0//fIIsxz0HphrnuB2G+pB4pR1QeP0xmdPzIdHbMBI2XIkjZDuJDsm32TQX5p0D4mqLK4uHcQUay
eGnZLirwva+gEPaRHnUJRl236vjoE4Qz18GVCKCrz4NxVdMBGS5Q3FUzQWh57PRmMMYFWA02OTLT
gXSQ2XHukvc2NN8A0t+gMurfCLCYVFhFLOe4vIb1cwoYA9nzcZihP9Jx2enNAr1G+j4VPMwTfmxR
QcAqzvuBD+fwb/3A2LP/MFNV6rCdyOYLPGtwp2UDRtuy50xuuzmtTXfzqABa2TGNWwaY7QUy0uz+
GtfrwozbJd1cxNfSchtyAHa2TTcJ73C0XBXHMzxBoRN7KRsk1EgEMbYyftGQraKuXxQADRxE3ieg
XJNLmJ4Qn89yICVabuTZ6CcOflRcxV+0AoeggX45eShU/lFRgtBGG5ycFbwMrhkTDck6aLQd1ppp
MjTJmhp7gLRa3FJbDWcJACk4o8kb6B8fLNcsZjwMr6n9XD2upJQnV8vycISkx8fBhHqFtIqmc5US
sjfPdp09tXoi1Vt75pBtNoOJbxR/WXH49SGIb5jfqNXypVQlR3itQlY7xjoXl4TaPEMFbIkYcHY+
mrXZY+v4le+qpeAhiwTSyMwvX1ZE3fnSYyIi0QC6aR97QioKDJqHiEdUC/nWloI4Qkpyo8nEMtwn
9sbGs0l3IQ6KuorU5q+WZH2c/tCQPoFGFpg67yGkcckHMQ/fZ/UDMLx9HBviEmBA6MUI6USWkNIh
mHoo3t3u51/0f4/hRlEjUCGNzcpKPRe/oP5juJFEHy1FSDKJIkzc0OVU8u6ciZVXjGKeXVEacP30
FKNuErIUn9OsXGR+qOUXKqjbpM49yJORVRoK6O/L59/Q3jUqxdeCrDXU0zrPu6bsLGNHmjLFb75v
OAnjWQ/cYf8DRbsbVdA6PI8io4nlwp8r67ETSqX3lUolcNOx4cvy0V0hbczYIIvnZKZzUCJ5DYwK
ihDRcUvzqi3eCpuNYjus5WqlrbEE9pAtNfTz/HzdAnvBRHAqlLnJUQXYcfjegjPP6muEsppgJVaT
gP1cmUtAtrg4BWz/9UnEUKlfzyWxX7eVPsdzewntrInI5Ct55bWdxBHsBIA+RKb0Pynpj4lrrSrx
sMD+A4ch0JDCtyVKNKTZKvueNDVpJPz8KJpDs15VNKtNMS/KBMQjebom9szjhglHOJO2RO9c+3pM
FrDaR+ipfs01Cz1NLStG6VUyUzWnX/uqAj55KEemNgKJgVKcL3IlNe+w0h2dmgeEjuc54VTVLLT6
auQ2BA2sfOkXHs+68OW8tk3eNUrKA69+HycvOXVapf9BWMMsqw718GWOSoQL3L8BuwyOpSGqEKc7
vPHeGulEP0mt4tnxhj/S+xL+dfGc+1noYIbT8vkc3IGVPkapKwRMId+5qhwm4c7OzHEz5zYhpwjp
tCdtsUnxGhAzaVdB/hCuuZQbvO6ssyApM1uLOKlBxhEnbuS+JQx7olcOFy1hnQRi8XxKbsKdv5Dg
zesNrZphkdYdla8MeTdTcbwMDCpEbbW/+VpVS7IaFhSuvSeocdfwQmI3yY1eXT7YSakGM1IgbKLr
TLsssQfR6lXlJ5o9DjGqczsr7KSnQiiIX0KI2VC5D3qVVZJkIY2XQ27pTH22zUFCKcXPKiFhNcY+
d7Xcjy34BUdtMAU94ei2pMlSzQGG/qaq1Y81gtgVMhyqNe6pJ2fDOocqG1hZ3BBN0sSMLyffPN9w
7OxN9tJyjVXo0+OI9Ni+a7YNtk19Z87NSsAi3Roe71A+ihQVxgyRHvTfELv69IQdjWd5FgFLb4Ly
sTDY0cAoCbbfooKgIQNCtLYqjwlRWTAM/QMdD2V90xAVOy7NgnR5/InC+ut0Wt4qocZEVZAvlmPU
S7jrTR22SVO8ZAQUBbK8nceXsCiak27wA5JwrhPiSf+a0vJq+0BWfW2vc4MZePhYxb2rx3kNXcru
/SpXnV2Q9l5H8dzBi2w2jnjpQrw2IG6X7nluDXVKQ7SZxgwz14DfcdsUnXDQZamS+3a7Ob1zr3Bd
JOHhjlmqNyh3ZcLTLwMxF17FMxrlpAOlFRBhbTDsjmGzcTI92d49R+fhWELx/9BtgbibGih/32XJ
thZwtiQGEqM6MCK2Y5ipygSbk0M7xBMrGwTC/MLYJ3eRbyasaArpTif9bJE0pK2ycG2/xcCpBm8k
odoJ+pHje/mWYVGN7WZThQ1euR0fo+XTp+aAnBtL8m94JPYwYzpmQNeV2db1L7F6nd4TboS1OAai
T6/7n/vSP5GwVk7DZ8emRE06284FMZOzWlyxNw6vE3f4YEyqbSVL7zZaoQhYgPlwSngCoFaOQXq3
Cql2bKJPoX0eRwuX7NyH4Vc2qHC/XVLgXDKpXL27QWnUh3tT+TQxdqRwWokZgOTWrHqQuXUXAw4c
lagoIqEno91Cgo1URsaBKEnOD2LnvSBSf65HAtVllnpv7YSH6m5v/xB4v6saFRenqYF0x38ctMiJ
/l/7VY/lfv/6v2Puo0oWLLhhBBJJLx9GC+/FikoRbnCqXXKZXYeSRV9lAATM8zky4Q23JN40jAOD
AkNtsK2ou7pitjqq3TjbXCjvg2AuSmnnZpe2YmL+taaQU1u7mnGGfN8oKVf7XmyaW57hqD1o2o3Z
0sxBULWQDIDGYSYpYQCS949btRxAHh7gFe3EXpYvgG79mQ7bPL3X3/cJGAuurskQ/AUhkxZkBKzQ
X7oAXX4HYF3oVx9OGC9rkM7duFohlY8flanls8Tk2b8Q8m+3fkE4bufv3/Hm/xByOWZtT6GAB1L0
AFUbH3bgxR5sW9CMCJSrBPSyHLX32d8th//vxINjNZAF23mMe0tHyqHZaQ+wHTMpZtldxI5MkNs7
VHDUgDn8fQmyhZwV4EXox160aLi2i055AJr2IOz8Q1keZ1AVn0VLsh7ehK6fWwl/2x35Mam8Yxyy
B7Nyo7PjWzcnN/uw8thh3MkLRvheDgzEkhKOHOD4sFCu6Uh/N89+b5c/Udv4q9Rk2HdJE1IhDX2A
urukNLPep33cGRfSwevS+BYhrCxNpNtIjgpY2fbfezJNFhn1hbtYgeHRBy1to8odmdM38Ez4KfpA
7TFxkvtA8hq8BuuxD1tK1Y+7jfaxWVG4+8VFskqXMS4ttgvAIdyZRLacil9eM1QkCkpoepi3253j
Wp/rx1cyr9ciHu6n4IUzT6RpZCdDUQHHg1yfglGyEfQHVhf+sPQkvzuD84Yglv6/C8jUrQV97Dg9
F/PjVe60E439yf62OnGVJXPiQGJlz/0HjfagbKC/G8XgacUeWFmsSPDiiIhFfT/gP8LetYPaAfEz
2nGk7u08PxX3sZODunPaFw/Ly2wZmzaB1+BXSPxGLUTRyHzwBkFN/fVRsS43iB/OzEu2XZlFa1vB
uUb/lMOOSbFlBKqfDtLp3qvDm1sIeYKYGbzDX0e97FR0cy5HlvcD4htpoTgikK4AI94NWWlRGn/K
1ed8qQOJaogvwQ9Xp66bsuXCi7vThBG5afGkAT+/80Ah+BYcRnvk6dizKRouXy94XhG2ucaiVtM6
KiuGE35hej/QIqHGCGM+TJBOb3vTR3rpXghtENTLQDEHNWLZnslMxvlVuiV9f+xcxReXx1dkZJge
u2e9QUphYYVUXH3v8qoNYwwJUxnSv/OAkxZD0OSUhisX/BzQLzRtakK8qcgp+jglpf3nojE6auIi
tCOPP6Redw0bWP3UveyUIiO3OqhaN6LGfk5frOlWyPoHlrc+A1RZ1i/NCTKnJweqm1tQQBCz2QL0
3grGgoSOnmw5RRiOvAECwWCjXavmNwPpLo73yBzsw6aMFlYavhD5cxoVIVKOYpC4j3dffTVeGe08
4Ij2Gf11DW/57iEHPYa0xeJwj3NOgHCoKfMIsZTwFyjk2UdSzAjaDfXVvVcH59GS/OYpbxR/EyhH
z/5vS2YbLXUboVP16XoV3ptBmlYrLzEYsJ7lBweBrlR/FCR2a8NjTeSdWmAgfZ407RDQ7FfIKDvD
B5F3Xr/PXJFhg1FnWAcqFfbBGvSbOguvNImIBSI/nLnoJPm8pSX0+VrRRRk2HXPJmgwOm/M82w0S
A9yGY8Nvbuut5Ns9tdmC0VN7CLZR9nh1Zmet0uzrpvfDtPT4ULTHc5NCeHgT4+IcN7NjHtbQ82Ag
KdCXbNHNOLg9gQwlT9caTGMvEAZJ8c/pMeDF2wi2V7yJkYkGh5yRtXl7REEasPvmDyGS0lno5YFi
X7dHfCetrGNWMoyFefTIlSsF/49VHHlz1r8vp6Zh6I3e+eJa9iArRU3SZ5WaNgDmc+e2lmebR+Cb
A5/j7SFCR04P0zsYSQzeO+SDTo5T5Gz6O/Au9ctS1eECIDmKHdWqXgX5y1nC09nCZD/rZ9eTjq7h
oUQYkZieE0IggmmYG4aKZuI7wzC22JPtsQtcR7VTPvuXD1wj+nqmJKhiuRvthGmvIe4tVDFkO8Ur
Kp3lHtfhGE7MZZORkEnf9ZKvD7okZRO0lGmQbgozpDyJxXLeUPxJGGhtpFLG3oIAfhaVN3HpUAPa
G6lS7FIOBfZvDYQjBfknshYxPcKhU0lkTNJPJWRr0sIycyBz4TTagDBWVxOCHmPkNKXBVHAdW0dK
IymhwXasXZ7oxFV2UQuBLcMtWKBpMuQ0OQ8nvFsyF+m8uTNstSvjdJhDWB0ZZvXxz/XLupQPEUGT
jBoB4lh8kSLljMSbkuG52t/8bYbhESuCrfJt7PfcRdrFIYv017DzBu/aN8jy8Wawi3Sz38v8eY4j
yGYsE6X5mx+lj4zErGKsoLsopuUheFlmB+tXGK4e33TTnPpsAsVTSmHc1R2Joj2TSkXFpLgPNFlf
SvB2c7HsPaWSXHjrIdXg/glk/VERs0y4h4fzGJGEo45YP4K14iD7yjLhk+BJYRN4JHIwSmZ63sFs
7IcqdR7XZsVWjpKfiGSHwE3ULEM7gt7rCGnE9I184tvVIT3JPxQ8v6a2dIhybQHczqWPKrkqA2OS
+ySGOTWjsVp8Kq/EPMih595FbotwqSsrV3Abjhj6tErgvRKNy4Rk0Ck49YDoa3oYE/hABdtNNbLw
InUGvofuEU19T38LLP9yfRQ3IB6oUwIqBPjvsPiBYrTATW5X1d06ObI7Q6Js+GOIP1SxI8nuvQRn
0OD3M54Id7IFYls8gE7g8l69O0X7/4bODdCQAWwUksLWWAK8wkghAJAXEYsaamd0K/Imu1S5BFqd
Iv7UPLWRaZCl8hYisVW7TKaQZvd4P8l9Nh5+BG8UsPvtk9kXVAc7za8z7ZbyP8DtQa4+7Y67trhJ
vab6J6cNsMxLvhDH+9hagQBS0xhhTGjO1bm6WC+wO/FouS/gO6WUhk2ap8wkTDAfkInreFzUj9Dc
wCPH+LQdJG42f7CQdv2WeOXZ27Aew2Oooo/7oj4BVzZyFEngtpref8+ckDepbssPdYG3yTMueQMU
QjbXoQANNXgf3ghAQPzn9azpV48n0WOux+QUyU05WK2ca5q7tmZkxH2L7+pULui/vfxTElbEHOe/
N5Fqg3VVlBgnsj/HgPcjdJ3P3IHlK1/TWvozcwgd8AKJoV1e5/Nx/4f74HMRD489y/xwEeWgUTmL
DZG/vm/6ysv46kiW/zrbTOz4UtZX1MOvJuNiAgvdRl7gLEole9UHENheJCwt7eSDIl0gdqdZ+JZQ
NRJiSXqDpx28QnvrPsokwwbhqy6H3H2gfArS3jrjoth0e1zNPhi1+oU+Im/4tEvbHusJ4V5e5AGK
zDxnJb5fY/OmJA5Oguh5Ij790JYhG9guYBg2T3EH4+/EKrRKW5UPerHzE2dhZMb4j1EikPViheNI
QyJ/09jQl9XWu+yGbYcIWF2Scq8kNmPC1MrWH3Xfe1JyHWBMKfgbA1SITYGS2XVvcRfQ3BWqswkF
DvlRwHE56v54EbXCdmMSMoBUBagnfSCopRuReMVRiIDf+YJ89Gv+LQtKtuB5wFVBVpX85UHb4irF
+qXd5FgfvVGAreHhQCBh2nz4tU6DLFUh/Da1Vz3TqYUAF/t4zMnaSJYmG5d+oUJSU3jBmyvUartE
HRkbtd/kP9KUsSm5XQNFRXYeDfl2CtZbiDKGr2IXnTF5Qe1G4dYGy4hqH3ezl/X6o2uAbX9a6Yv0
y9QFy9DLGE6CEo+SM/GzSofdtf+c0RdLMUlwcouPDus/M7bqUXUQnfZjxHqETEEZMQOySLlnKpQL
JnAsE7V0zoARIaYJaXt2E9E8pbljQKbc8omxf+HRmLGWi7nmwPevnhHpeKELnX8SUuD0N4V1ii1t
OJKjXqK/52L9el6ZB8NQEO8RLBN7rZcLeL2fRoR8ZFkxILF2wA+ZAgcaGFwtXtqXQvHnH/h3IbjB
s6M7w0Xk2CdfQz7LO1lFnVT5a2DBH7W5dd3FXWapz5TYSM2is+37E0eL5JfjDUvWwTWECvX5eaqo
1IBjHkhdl++idE7D/CJELswuc39IAdBk3S2giS8kXqR3QuSCU3Lx5A4e14XPefKCVfQFwaWGiJzH
IlyVwEJ2a2w6f6+/ubpWGOsPOi/Iv0vr3FPqj77rLRPIhrlVp6J7IDgNWSYcKl0sCRp6QJRWy5f5
lOZ9MDj08jAYou56WGGN+5fgbbsTT982eI8pIJBCop5HUWbUuF0BWcrEVbM0Td2dCYaBqcbAL8a4
pgy02Asv7v7WLSsSC6tXTfvZ/sG6OZeC86AUZFWP98WhPuZW9vMU59Ygi9LUQddhWqjlJar78FEI
/EZ9vCS/+4IX23jMiDm2Ac5BNdjFbGxij3gR8LTXL8g03/ZsgUKStXoGgbHO5rQtJ3b2y5iH3sXl
0y84AeDBYFV1m9ZjSCu65339pfMlPqNlStWDZ2pR4H9+P2jQm+xo+1cn4VlhZTZF76yZxSOIe8xb
PItzTm/+5XSoHhH/HcfCYdgxxvqr0NuV7YGgvC5aNWi9R4YVnPfOZGsCrguN6b6+5Ni/EuRv2lHg
twECMVGDXTMSLgaA/XUw7p7hyGtSrkkMzhX6E9vIEKXnG7u7ohKQKHTMSl2beBOEMeWKZPbN5JLS
bV2QktYERNzP06SGPJEU3aHr9nAnf17hGZ3T/HWIqfjrMRlOdy+a4fgxVHM6Avx2lvNHEeKpKhO+
qyLyM5gxrdjMRrZ3P6snnw9Jp5r20mP/c/PBVVZldw5Fd3vMWtBu5as0bJitP+vTxpGy/zxgE/oa
y/iNHYOFZt1Va8+YWjJ8MGJ93lbu0Fm69avirpJK8ZnhOqeaM4uUZby0wuAKSYj//BT/xcCXLgnA
s0RS5BU+tDcvWEdRRPM/UFYr1C28S/Enx58RZM1Devn3xfFXTl50+E0N82JgHYgKzAVNKkZcvBeH
hwUip/gwi5Qa7Pqh/GyvYn4dmcw5/1oJQZ+yDimBbf9MuaR/vhJ7DdzKTaarki8qy7/6AFrjZMf/
kUPUWIkTs0ksJpLtQMEMfVKGiBH5dBBwUJdoZZxwrS7V+CruknFunMn+c4oAbf2tbiEkO8V5CN4S
4xeQDfZ0q4PrNz6v9niY/w5V5TKuuYpv+zcXjDZ3DuCdqMumh8/CJXjoHLU1GvYx82Qf4iEyJ8cX
g9FaJGxwnvbRFOBDu/vJCHLOEwvs5oNtdzeo48uw4j6vUlvEEMQOCj+pp8Z9lj1FDeQqqTAC5R3F
JAFm8a0JYMbvfVK7FpmWsiYFSflgEPkto7V1L8ypaOCXi7zI0y39EJytcq2Q2lmdAyIsHC3hozyO
mCyKx12bJf7OHwnJlOcGI80aEZtmelEYmBH2TKgsc2YzkMnp+OdIbEHOVpk/7AJynQFjjcGct6Y4
XF/bfr4rFrSXrtPR3f1jRtA6hgJRxvdhJaIQBf0X5uBm5C0WhHFdjegsVPriwSt9l1G99Ybe4wyP
vgYi+QTG+AY6hVA6B7vbMIhB8lkS7gKoinjmFOIknbEuyCYrNutijBuKj+Q8bMDUqInsiWwWVkKc
7l5nNDDsTlH0tiyITj4bWef5LZAB5wU3ZOAf7Zd+jTX72+lldpWqDtBJiwH6tHXrLVMrEGLlq6D+
GRPcMYeXRJOSmCWPkAcVQN3jfPUEHCAC4StCk0xohAPOmh72v8zlJaSGwTfyY8BBz2fPN/n5BeyW
bOgb686618Pt1oh8HAbuzAoI+TszUqMc1Yw2qFy40zjD8v41dFoisZ9f6IfT/IMmA4xufjWH4yJP
AP3Sgx+dZaYwUqGfd1Iyk0LfqB8SxFfvhmPr6smbvzAi2ahLd/DJh581ayZ4p7It1+CxYSjLFbho
XGjbXgg+9S60k7yCnX7uJivYbY/Jkbw9jUwr8xzD+SsbLpPOTIA9bHe+0ljiEhFzEjPMDO9WftLv
wR+9UrYNyxaJpZlFiTHWW+lFRczo8MVAdFhTTn5D5VCfihwsMIOW3Z1+BI3oqzZWxRT3YOWrTB0Z
jkJgn+w7r9XCdK+Tx5W922MYFqe27xFaAwWNpPbNxz7p4ModB9Pc4uo15IVE3Y+sWoxGODLjleKv
IYbNPDFmTq8pt2mW5vT9P01qCOIYrc7/cEw+e9Tidh82aCWRus0k2nNbrQb4rlt9d2wbexvWlvp7
Y3Qub0Hwx4+Mb5lbXKCbV9vmgH2QraMkXlkZkwLsqb+X3Sqt9LTaYuQXg9xKBMn22Z+zc8KuMSWM
dDMiSMz5m78k8RAl6ihsg+uZzexEcwAxcf+tFeGmVFVKRMFTvymWKDcDmqwCrv+ZbVVKTUvRhKMS
Yd7zrRh1gI1dy1eyPMdhMmTPTsym2YzWygYDS/vH20ecKvJaY6fN5jZ0omqSViC0KTEb5vSdHJ43
4UNnTlQpAh6pCzcjDTEIUau7jh15PKbH0EYu82U0C6GdfxYvnT8tu1zwGhbwxYDN3pAEUBx73TSI
hoqhxccbKYvc0TLrcaGT5KcOC8bqdO1lxq1A7LiyU5UAY0AI4XJev+aeYWanPmlwhRCKHnZNzHhn
548u4PkZjZTrD8ArHszgCxQNXMhbvYCfyE7sECxYKRPWY9S7DT+Wzwn2L6lkzWZNFEXYpyxpgzaC
iWSOpvce9e3P0S3GmRofiQWDdBNnkPF7UoN7D+wn4m3uKFWTAS03QABaUC4DUffxg4J9ecWdsn2c
QYUTYdxjpZz1AS/k7ByFX1bVOGMhJsedHWTgBYjemiI+V6cDCef92E6zaTy4/cjf/V1bYDIib7TC
Jg4QvwXcgfqwwJHZBiI1WWBNALrXFHlYsP0gLaWkG0102ZxumblXdG3a0J+/npJ1/WxGmbXqDJ3f
VQurnKcWPZ/G4UYRrOOY/mWhzSqEs09/7JWbSdjHkA7AJ4j7+YE8Tdhvv8fTzaHVTkQwscvNf7UZ
8TcRvfuSD8AZNgoQz8IG7TxMstruHh2GFhB6JLGgX/XC+gpVVh/9GbhATXKFsHxLaAJdiAu2nMjD
m7sb0sw0levL3fhqOPYZaEdikPpPubG/PTqXljUw/sheVAHJ3SdhEJBir+jDfwvReCAy7V/guh/v
XssjTsdZGxzoBqxtHcWEcW/G9IXMd60RZL2iVydg3PVVOdIc5kpZIyF6NkDkzCjBN92rPlOJuB6O
aez4K8Zz6CoMsSRmlbRh/qnkCMVbzYDYZAFBK7ixo+4NPukl3BOqhyFVEGqvpeouyLEBWHlEWbqJ
vHLIcUcOrcu+/vNqo5PofY6/aJi6gm+F+Ef8qaa+NUZ7HpKmc9QF1+SVUxwk4uquheSQipbtBGxv
sJN1gvgad7W7EiNs/2xaIr3VQAvmx+1D/y4TyES7FR1juUFQ82nwEHeleaSRO+2plG0QK5i84oPA
fAx6kRrSOrd5MHbYqArrIGLiTHFqsOAb0CMn9eTLpZR6YYM0da1E5nGrbe0EEAaiuAr5rOL51YzA
2wLK0aRmrACRNPMQrYALc2N8KVarIPONbZ66scH9tqqdXeZOy8AXOmpm1ajJbLehGPQL7Mvh5Rnr
HIY5uio+wM+8TWUAQKcT86xBb2TLjSU7+FLPPCkmUnS2fWKThBTmSgE5iHXuAnTZkQ1OHwcBFBUI
ua5porkarVe0L+ddt+h3PIwpy7v/Dupj7hm65jZoon8mmithPchHXxCQyuZTK7BwJx6VeGZk3XV6
bN5nSWRkeEtpeoOYjekKLiUVpR0DF9M+OCxQh2LC4DS2e3aLhUHRjPBLOqRiTbsOL6C68POhCXf2
2aQhvPpkbw253+0b+yM0UNhNCXQ9h3v5aHFUP2GNY2yI1V0caZ/6iIxSLq1Y37+vjYCWj4PGavnM
wE8/ht/fgmlSgSiObU6NQtT4qe7hyBDTVQb4FurC05eaVKpv0brgfiwI+2bhEIfwtMppqMOG+R6I
mFWzxvJJkupmuHwiY48nbZP3aOFRGFgKwgZu0mfXUO7UQs5Atc8TQ6hEPJRpMWpU1rw89zLiA30O
hexa5f/5gCrai40/WO+lft2H8E3nxsdGoIAwxxKtQrYfBr5oo/adSUpLxOP2DpSe9slQGnZ8Qkx7
PhZ14iZ72Uj8wzc4FdfYAth2ALLkjk4GxEKedFl4VzfynZxS2Rgwh7M4jNlK/3KvGt7XJvJJOBi6
KGvEEUdIluzFVDtRkRSDIQUQlQjwBradwyAEtpZ+0IfEW5cY1Ib3KOYDAadYmer4qgUizpXRsEhU
A+Q1NyQN8hAsNfdK12Ew4ebDKA5Pf9E4PQOmDOs6LUZ/VsJmXDLhQqjeC3krHbI1CaH1C8CVSfrE
MtwfVWmixZGmtJovIbg1UsZCwjKddEw00rPx8C+ceELWFWEP1RyZKncE6/kCm6jamDBBApYIoxpP
CeGsH8ERNTwrMykicBEGB9xndjZ/jY1NUXdImfeZPSUJLHNNL46qzNDJGFmIksNqTrSpI5lGVziO
fqYVI1PvRw+Rzy3Gl99fWt4m16iINjZ38q13CxynftTraWtQ6CARPVZjA/x2tPKc2n62lcIlPD35
aQJasmy6nInE4q+4bxNJEpWOZM1Cn0orYEYczzu/yr9EhrFH5Xgw40aZny0i8wLkr+eXtJfigvvq
qpE4jVFgYiy/I3sN3Q8137dHyS2GXXYEXvfu4AyXZaEzz3GsToYIf0achUTPicS/BnbNWPwIOglg
jriFAN/6ENm1Rogv9udQl1FHVn0MMkaBV7IsQPIHZ8QRrCGs3CKvRCLV2CBmmpjBgO6KF1kSJL8R
SZczTHGVbiGaSIqdYbuDAgoC4+sK8hWCFgJZzKbFmRXpaJb4xkhZ/Veq+ZOxdxd+d/KBFPSskspJ
0+S1ZX4/9UnDouiQCqD0q4FSKR3MpTSgX8BOT0RP1F7VpbQNPjeYOCMO9CXQn4Hl9N+8fvy0vcK3
pk8jLsZwovOUNBRqCQXGQlpgW6pzgLaE4Sy+ayHBg5IWcowN2e2qnEB4V0u1qKZQCrCvJO1H9NNe
/cFRtPl3UQNGwnmtdWqKPmmmrVhFKBoJKcACN7f5vziFZCNF8kRBbqBp20WGRFFEgSdRP7atR3xl
vt1+OkCibCNsHBS9mMvM8OO5tIhEwfobVa8Si3kE5Gfp8VJX4ASgSOrVQzL3kkAUuu69jCokXpwL
mgs8sHllOnWx129tKTrbvWnBZ4U5tGNtTiVPChopwH1rNOVSw++10nzu5/BF5nVht7aCuAojB+Wt
trZ6cGARs3BvfiPEOVLvn8fN1qTDuI4NksRv2kRObyUZe2Fy6uWM9aH+9ZjccNDtlpswYS+d5sq/
sOFaPfigL8fvwnltZvPDr+VwTy/gdRL+OvKAJVxSBua/WqjuCAtPouyYMY98yF3RAEHG5bdPC2K/
ss4M7mPTkFOd/wd4dzmdrwgMKD9SLzIBQLdkTZJ7whwO/64LmmvexutGOkeihEmItMNf/qwlSsYl
k3Hs+wcyjIea/aOkUS4e1Pbv68lYkKP2sODiV0vD9US9645zB2c9MO6QfoSzWuqQALHdZykkAEtt
4Wr42fao4b5OdOps7Sk/HnqGGhDfczEVVkMal2SX+Rnjh7m+mH3zv4MGrVWk4SdHSXWPr1xmb8eC
5oZZ/t++Oe2sZYJlAa91iyZhDyLof9ZeFr6LDzkQUozzCgnVqAvebbZdGq5hKRdTsdC3q4aeqnGp
V/h2q62jZJYWhbL92RJg6KL/Ka1yUSwKRwOjkph/3xFUMeDY0e5Y6/88GxJPQb7BwAhDeL+exedZ
zOR8ZxGjrr8Q8SktbZiVCxsEDHX9vudtb95zrFQ43f0ckf0cyyJqN6ZDR5xLJj2POKRYFgfY8v6l
O29sG/r2m0C4s0bJWnMtMU+jUnOF7jY1hKBX8wz5awo6ZTl/wxsN5WRlN+4RVIp38GTSJ/91AIOE
YpxJNgdOOV646jNGrnl9d7vs1aBAz82xX+VnBaoq2m99sO//c04+VmFDAW4laIzWeSnOoc0/ZTEo
U9AAvrkt1oBecKjAZz2wedQUJ13GDupWMYD6jDxOthnHl5VGAXazrOsvPDF2gNQlCN26gXunL7wd
BWF0JcU5rPMset1mWT5VhEx3Kv35SBYwD3O5AfrKgq2OAyG15zt3M88qCwjG2ysqrxU4i/J63XwJ
HEAlIgE30W9bQqr/9CfKBfJWw4evM5uJ8CpBf8jezuvKXoCb1w25IO5B3HkT7pMPCQZObWAqaL0F
CpxySt0LzVfUjN1k4hI8wOCWvKuIbT7txWMPVfibpf1XOfaHprv0/XT8rD/zGteokX7G3Tsxqqzr
jQPYtzE0rhoEjHE4r5r2UIpB81GEwvLRbxNMI1jMPZc9mXoRY7Lzs4y6nVG6fsiwUajhhZmnKSnE
FWqCw7JtIBjCqaJICRwAfYULmyFd5lHrDbfzPDRYfHZqrJyOCIDYC+SsoDwhp2QGZrtjZuA1oNme
khyRTeeSBtS2k3Iug5Xhgv0ITkG43qiER2VdF31D6h5TM+/KFsk2IrE30Hfan6r75WXN8PvOKHfw
lGPJHZ/4HvHjNXGjh9tvn862ipVFGYRZ1PsfFbrlBoLIUcBLsPUjbQogXFNFFQ16AJ0dWqZ4IbQ7
74lmQ7K5U3T4VJBxAeT0WiexN8zp5d3lB7BTNUpGB6JQ3T0gPEZyjJ4NTSTr0IQn8eNwxGtTrXfx
pxGl8VMZ1grnBHLG+JZKiuKbHxtVxv0KGAh6IhF/vHW7G8EEuHlusC9l5x3tocWyVFKpH7JycaqL
f92b2OrcY6DlHVD7mwUEKLCFDWiH/7JUoSREf0vz4zgRdRoQaOw8SQ7QWoAvrodOFy7BnxaL7vSy
MD/zhFjT0J4PURQci3A9APPgaAjSn6fKK/7ofN5X/ko0wM9Fwtayj4u0Bx1fY8TRk26Zo93A/s1H
V6F3OIH1Hq9Xyovlh9eAGkwumBuqa+2RDBjCAZS5a4cQM9fyP31Y1ZZ436RH6/FAZDekO6wuvyJH
6rbOyOtZuF/+YlDclNE0ubikpyBGMxK7Ic+tSWXnFzJxPjd+S7IKtHi/oPOuDBbz2I6zEcF7mSDK
NRNMyLADycF5FiGJn+nFOTZbp7EHe5sevpHGtepJiCA78kTDQqzXgt33KgR5YrbWrdPTHzfu6UVC
auc/gnM+iVhSZXSAi12/4rKpU+H6kiuoTGu+BrbaIWj4hO3AuGtIFBln6BYsimkcOcR5vHIBnCqn
8wary4JuzHdvG7pNHr9J+lrFfEACxzeAtWoXK98qfZUr/SZh1mdSkZ6TU1B9XvbB2kO9t0lg8FxT
IeFKHVmZgn95YYMS5H+gNgPU4J3pG+1rk7x7GFi/BQ/0cNYql2QH3eHqV8jgcolKRNRs0mHsvWXA
xTRgKQDnqMtH2N+S/ZAZ8piFgtfypBruObgXHrfABTgf/Fd8NRzWMhcLMnI+krBByLHfEGrzrh8F
dFbFDJccIiaFkMZZCV7uUcST7vchTqTvMVem6gPyZQqrb+kY+xfbryUGLIr4Xr1EzAkHMwweC2LO
36GuSMa8QlmhMHhlhV+DvJ65SmvhPbQWiM6oYL+9/9jax90HvrKGPFF6gW1tp8Mfu1JMQkcp7iYb
tAlAlBYpQAgvvN4v096YcE5UJW0qDQx/HeW0h+U3lz/mDTvVQzZYn8bPB+Q2+71h8ug5QRmuqtHi
5jw13w1IaTlC2Jgk7lUxqgC9CffLcNjLB5A+goqGYeEZ++QUSQwbaYr+4OlNRINXdUq8m8chHLk7
ehrwCjdQpIK2AUm0V5Omkf+aVBIZcoCUFi1UOD6KuTlubu7IjeeyPos3L4JfkpvtPBVkRYce7wJ1
GzeNI5TFhG6ImmoBUXEyFo6brH9cR48qYT+BfpeLaRUxu81t61RsAAfN3lat6SMUav2UacyJfdwA
CSzFasaGXCJ6ExVI4dWjmF71PmHArCT39UeHOsTrWhgnY6NJF63GSrkhjzn5bsuc5f+n7utKl/o9
uGLofgLGqDfUutZOnBO2GSE7DB0uAXIyB3tUAAASuyCcT79fkQMNcA1ATmU2LIShtBpidJqVbNPO
Cs8K6/r3neMlcm0W0F7JMXVqYVz77u2OUZWun/hVDK6O8T6+u+64yaXnwyLvPQc9io6wO9n1078J
7xfZRA0hfTGq640RzD32xxJu/e2TjOGnLGxPZVWrT45b5Gd+CJdFPKDYeejNYQfc0/AhrN6AJsUf
djmW3wObovg041YSU8p0Z2L+t+iuYMr+ewCCN6rDrjXgEt0plLXPAOuJveSsmqqk3RMGj1EoapaL
QUvaADtI3b4ExRGSCVSTx0GekCSYlZK1bYJQr7aRmnvlioXBqod85+X6wbE5qQGFU+C8G5m/ZVaB
4yRBFnDSEYs58QGLG7YtNLgqAQEhBksyLo7agF2Y1Pm0fza5CK8RfxTgcGVBMdQB667JWUic3uXS
ZYfAl6LunkwdgOv1NtsyERLwZ5apD3Ht7vilebQS/iWKD9TDdG4bkLbLuyJvATB9xBIj9a4ebiOy
rTUPLCofz0eb/OpJFzQhJRdo06HAL/En2h0dv5BHBAT0dcww3H5/LWt+8btInDzMtwVni2rF0mfA
+4MZVXpsvxBD5wTY5KXRgprxtjwbCjvgqWJ5A9XMZ53HL6Qj84pRvOdACUkDzacXpzMwYjtS4DIQ
n3nfrZH2vOAchvK11X2+SRSnbXDREvtqZVPXTBn3a4KVQrk+i4L1Zk6u9oS4dq4U6SPgvKk3wJhW
BGvVj/v/2df4bI1CjYWFVNhl8FmPsuMXlrSgpfs8HHwtTr7rmArvenh4Brnbm3Ig3xiiE/GtcK/+
/egM37g7ddNwpWD1U1FlGQHedRPm0HMi79a5WUSjKrxFuRc4qLutaznMORiSko8XtsuCqcL0Qt5p
83OQopYWroXfk7PUxtIjvW5zuoCB5u6VQvn2MALB+SRMq6rvGj282ZTzkcPoXhdmMVnruuJuBGoa
AJP81q0qJSCv6XrHSsfN9ilmAv0PF5ViIA8fcs6DJ7/Wu+x82zvaZsLmgnKCHjeKTVCQ2N/8rl2p
Uk77b2Yj1CKEFjdxAJ8GyJzMYCbsFa7i0LX7DgGWR8RuY1u2MvxcSw/meXYSFR8N+HyUH9aGkSlq
UWPmn8jJf5KiKXpBfvBtiNZSBbtCxMJPaIM53+baFIvsL3esmqB61RS+n8IT3N+GbNA+azmPgSa5
kxHbXhVvgessRo8ik873m+XU9ordxV7UTziPZXL7aTDaw/mT9ROhYnZtyumRU4y5LJ8NHo9HyYF4
H3XOHu7M074rrHBa7kavs4r8KJAEhkVtDVIICUfxfM/w29SdOpj/IjB9+Soe82YxfSui95PZljTf
IftdaVIvXLGLRhrqEcyVRoPVoKvopk7bOcU+C9A6zq5tlT2i95O6ARV/gBI420rx/FZZbckuFNX6
ScrK/uohWHYp3FHYaMNbEs+T/+L9wwG2j2IzWVj3mG5fOtSCeVg65JQdTNPSUI+KMPahEbXfcAO9
Jv+QBkWOJRXxuk240PFnahCHp1j8pPPl5HSj5VxJUzb2RSUAInyssaoQjeRBDjriUVMPQvhNg6sO
JWAlHfbF8d4EuvJyejNzUZow3j4bAxj1njT63/TRygiYNHaOG+kL8pY41u2Sn+RpDub0QCGLqFgA
MdT0Cho65meqZTosjozlJUuEtozbVmt5PYX5+k67uL5joNv8xsmOFXwgzikdZx8ZSejm2lz5YnXZ
u2VM/iB82DQInIYUqX0/5354UxYQjGIVM24h2sNu6doaLSySM2v4v6LnahwKX/Ix4Z/35Gxv4UxW
JjW/JeYHK+ojNvqQ2rRrJDai5plga0cDdgn1P1edugB1rc0eraflpTaTnKwybcq4EJRcf0p7dB48
xJ7ajcouXzlaZUFUoDHUhG0opKY+bImc9jnrvzT/89XqxSk+L/j7Ms9nvdHpWMGCQ0ci2BfQTLQY
fX2jn8TD6tOMNSMq+oJVqUpGqdHn9ikBuMu5IlrK1j8OToj0xr8giMpQ1DhfuKEGDlxkwcyqZLIL
3shbzNiHb0tWAvnEexJAVrXuImldK4e2478LkQBIyw1PpchcecnZ3jBwb7T4CLMBBjjNm2Ibna4u
gyoxqj6H4Y4XKS6xmsCrGxmzeNcBU7MMZpxSom6IK7UrIYTzOSeI81bB1+0ZdbI542SvfY78WzAJ
XO2YFtsS9hCcJICt2nxw/pTJvOiU1Ie6GTrLmwfqieomx+S/XplP3rSrlumIa7/J9TI49mcZsT1Q
yoGkp90dqobxS3RRDj9wuMYauAvHmXPiE6r8HM03pbSvQQjsT2RdnfoAZwwrNf5I88nC3S9I9nPO
tvBkxp1rLB0FbBjg8zN8SSEcR2O8Yb/lheK9QjCP9XzRJjnMlYOwkOmazfObMZHR/vXpuAb1FIYE
KhmYMjezIUJ5AsSMAl+VZejsW9pqJcHi8fJgGBIbge3QkM9a8rV4TLJj/98yv/vLeTshZwy7ZV8E
bWgXM6qSvfPDUKKPr9iGHDjIhPP3ij0u3HARer5pLU3K5UCAzZQDiAI/EKspwYlhDc0t0P1vXY84
4muheSo1JEDhnIPZ+qo8WRWMWfjpfZrCczu1WbKM1rlzBPJtImK0vzlYHbod1e3JA7Guhe3kzM8b
BgiX9LUsh37Po5MoIZRFA9i2MTN1uZk7fwaPF6+d9puIzNLCMAkW6u09jaTE+bIWpXYlpB8ma8cx
myxRVRLTHIc/Sr3BgYTJ6mYPZ2L0Dn2fkfERyU0X3U6U381e8ml257HjWg8CNNXZw0zOBQywtA9+
LIzaQiB7Wj+WvCmipYh+dmTKW+RJHsvY4Zd8xAD3hiTFrn5pwc6oc6nt8GR3mmqi7c3KQUAxTONC
Ya/4rZHam3ZU2WBdKPOMCpUKrkV25NJ1IIvxeR6wIUY8abXft14HkFZFAkSW3VAwqpBlkg1VZqEt
0XEnwZt8xWjQiZy/kzXzARepr60iHVDTOVxciY8afqi82si02vBDoSJUD45xQG5JS6LHgr8AD4pL
dg/ZEFin5JtAF3ObMUxpi1835krNuk7qVcuSGtB7CGZqsnlRz7Emg8ljQqH0lUIAMMSn8a4fRHmx
cr2DsuoBRk3VeIWHNeAZt+eXUCSS1t8eIzsw2LQ7L+ys57JKfvyVKATFQDlo7/ZXZiuEU4JK2bLM
z3Wgps0IsGcxGTpxBmCeJe9p02mBSxXydPPPJ+gwWBSlf2gwOTxtqJzD4/JuVmrD+9zc69wiOFpa
vH9ZTrqvrpT/v1UPaMS9fmCzk92Nrueg39ku3yMI9+UrvAeM4gWcdy7w4ulzi6pk30wpOhfu5jVX
9lzyQg7SNxDRh0iC5sGTOOe+Vwd7U4H9VBSK24zyarOje1z55aZnBi35SmmOSqMNKSvHHwSKTYgT
hAX/aY5ObjH335oT4cLdGNEFEaqxPeaHvjtBm5zECcmNlwaQuMBOnlFA3kzPsY8FzT3CMyeOZNEn
WnIFzC5xQai67vv6MqhbQrLTwJADMPqOaqt4chYSp77FZmncGhxU9NZdhUxXAAMesm3XN/J3xFhQ
3DShAEHY1FZUCuZyzuu8mEM2pK70iGAp1jRKoTra2OXZhQWHDdPAo7jWAWGI3sAFwQhVX16gVOwm
uffA6te1ZmWfgbtzlbonoD3Z+yoEsX+3oGRFJxyFdW0bIg+KlileDs++POMYmlRBKV5jNKrncclK
JItb/JdP1cgMV48JfSATrGMDKNQG0OdkHydX+vkP8X6wt0rXN0sqQNRha1BgR3UO1cSHcm+zyE0k
Su0mBWY1SQbNhs4fPj7hlZ1L331rNkzIefTrXrUVKwOWQlOJvgZ0i2D4Q902QBw8F28BYXpwxJyT
DRI78ealFus1QOGhH002O/0qaM2g59TIGvSgJlTzIl9Q5vvyHJ94GpJ/M5QIZkcvAo/PNuhn/zg2
LRtxIyG/wGWUZsourbHaAKBeV9hH8JJVLAVcE5TFaNtPkDgQnDD2yFC2e+t5Sez4ZprheleTzdtN
69IiuT3f7iZxnQeRHtdqulrwIWw3/HwGH46qBGhvYg9TsQH+fdlm9TpcEh6ULcfoglV1qo84oC6q
GkQKltmhYPs8BoYVgXr89wwAuea4ZhtC7dXFO+mxzuv8xfFVwCBTvjj2Ynz0+9keTiq6zPhMQONk
jL+5C5FWsKL9Vq4IScLMiNbQadFbbHVCBFqp52qV62v9ys4JSOuphhF9DO+g1PHJJg2NDK+BWHje
QoBl8JJCB5s0mWDDmB0mevFIkwm9JLMkWIBhGHQtF9vl2W8uqslTqW5NrMdNR77S/PBLlNyAqPOJ
ji7Vuiq+oyPq/pjZ/LMlhu5lKleff/uTpnL38zaoy4rPF5SD3YkU/1RH7wi1oXxP+ifOvZTxl2od
W3k/6oYyYlskzSkyU4ruS4eYfMweMisifTrTYeZGlt74AGBQ1KbcjXtB/rZpC1zSJvX/Q2sxjZS6
eo5Q1E8RB565S47EmgctXqHFQRKHKxdXxfL/RhZyemcgef4QGQZNFbw7wELihkMcdtIqpPkvNKcW
eexoTrpmobta2OgBnXwwwOu0o1ojpWkwivgoOfIa3F/wHieodEPxuwcML1UZIXjXXInAmXUdD7wH
hktJFXMQ9ahP81EOe3mXn/9osGgPduZpFtGRhvdg/p+s+ZWqatSO02F1vI53MDjUhhrP+aCv40dx
S5NxxEgBw5m4cgIET/k3dVI1F+4AX04bi0VbgNc5DnYUS2oE8VUYaU/aAJqVLg7kF9zt2CO12E+j
lzmlk8dGcXggZeoFaNyHnsKIABdFXYXzvvILviuSJFUuCUkWVtfU2xf0Vh7qriQJJ4CI450+N+O9
M0+E83Rd34/TG+/BO7hUYY8ueMeWNRl7OFK6FBRaV5/EjyEOWJubGOQvsHv7OENaRjTPZ+J1GcyB
ItITT2KGClgeSe1lgoGtKj6BNnE3Tl7k/VbEuWOwKJxl56AKTQDd9A+UZElv/xNl6DhouX6zIfOT
EoSCKARHynU3YRP7CHAh1jlY951oITSUE0yx1cuE7GEh5VZtDOQojkp1t7B5TQdLYB0461GBkp4+
qBMyN8tehuwryoZxpxBP9CwP18XMPNHU3IwbXlKWbPwq3xaEVlFv6/5pZxw+rrGtSgyYUNsnUQJv
DXsRy1ZD96ecJnB6HiM2kQjuRhz0NwFqk+1sCsaNKxNSAYBeFcn7Z2xYESVssOaUb/8jrZTeJ/yE
gFpu0kUHw23DV4vukeGzU+fVMCzFYuOYCPZQQUfz1L5QdEL2S7BBGRdaNPyuBwnsZYO8smA4F7Cx
Hg3XNYHAynYtCbHkqBIFo+ek/zH2RjlPZxFpV+KhKAw8e0C59Y003MZh52PvHHmg78B5pkwialH6
/T1+iQ6Mnow9K7gbAmSnO7dh/5ggwt/CeEnWSDvOxq7bXhIdpwWDGffEQtezf85WlXJfxjWrNf2Q
ZykiqeNgc6wcxAFy9z4pR8sIf2Uucx+2I74kl2Du1AzKRWoGb85yh3b529NVQaWZ6/xVxsWSaAfh
54bXiUb9ZA9ThgoSwY6/5v6kgcoqfIoQuZV/wc2XKsbXjxVzUmrv/WrCddp2TDtpRDKBRpFKpILI
WHQK6mjxx1wESEKBQz/ah72A24lE5PTxWGNzy7sRtP/7bl0OTiUuluqx10WF7LKuoGLcVxjrgsRr
sSIEoNbMedfjIsosYxAhUO6oQ6r8fafGssI9/OaGxsoJ7ILot1wP7rnYdF3mzeC+r9STD4B5X51x
owErpdHI7vyjzScFcXqlwpIf8OA4hYJoSnt+quZ5JhrzIUIDsiq7bEUSlJrYfaOKeLxpWu0fmfen
njeCdHnZFBQR9A7V8H+xuk+7oHaAWVXP/QomKCV2gmz99VwytKJVSJLs+bmfxuLQTLX4C4D068uU
QUjUKa8rUzR5qlNAn+Rew8PQty4Lt6JlpWLuEeZuUNnpZOGmeYvypiknlb0wWJYaYOb85AjTux/y
Nc3FuK6zdXjCPn9sjANEUmbpNs8wwJKZc7Z7uiwahpZoyTtFK6sIDx/lGnQpTdx93FX2SUruJ3qC
oGEwNjq/mb9t8p3yiPofZrEdLHo+H7i86DZKK9CPH66tv9kS7+e49G/LsESwgWGFDgtV400N5ukA
n2ViY0sM4zTzOYZxZrh/TEhNjy97ccA5MfuMmUY4nfJ2zQpgjVEbY3fy/6JjvfH1n9WHUdSZ3qtp
IvDCTccsAfJ53lQ2Q4bJQi2dCScBcnCT5qnRaQn/pLICgiI7TeRrSySmok1mYe4OtERf+M43tplz
39YLpw2WwNSs/7j0JfoQZCzjvhiNJ0iGIDTvVsKKV/oKNPw6Is95iUVB1f9iRe3uPY5bZ9RN9WG/
PazWtytKwTISQTFC7KTFF+iliQct23UKQMMuoc8ZqtkdJEudNfYT8bGHTuhI7pEyVriqORuvphfa
4d0inOO39zTNAtwrTfIe4CJrDpC1KBirwyI8UJWiygeuwwZ1LhXaFmlyyXs8W3Ci6kzOPK5usPxS
t6vNLx5G4pDFaFG2iV+7/wRzPwJZXmpLXTAUDEd9Zgauo1lGAn7bf/qQOEG+0m2QFAkEpwTS9F0d
vUvFZ8UKn69YkrB48ZPxudSFhSOZakswQlYzAtwUxkA5FMDXg8GdSoPe2TNSkHhmG+wuBZVgzZVw
fTMCLpVpmC8rvSF3URDDs6iXUGyVwHlnswOs2Rxu7qgwgiJ6xUClQldALyAMWxTWxg2MmqYYCYvs
F/MUWRVhZZMIG4PuJ/Ekbi0eCpl4439kgDtMJn8txQH9951iQm9oADH2GMFTz9O1dW8lYnQjPRok
4+TW2vqfLo3uHr5xnN48zD3mnV1arLswcn5294uzkdCvxLMfJHgJID6DLmu53szbK1RCgqJeX6P4
WSR/+oR9D6M2d09HhuarW2eDyW+CeELgnu4zrShtvw5ASFuI1EKJTStrTiNkCDqyguXIXZTy++Y7
Cg11NY3ANBDxtQohGjOSWUX4Xowg2AZRDO6NGt97/kgMPI8LNMWhHCqIja75H0hPT03JqQv/UysJ
rC7bgqm53pwByMputWGn9pVYqfYp/TrmN62xQcxRBoLXG2k+n8I6lBoqsLRvYVbHWPp0ZhpUDDjb
6BUwIlx4v1MrFTUUq5kkZU4yAh2chjDkz5gwGT3oX8VudXAN93520747yhp/eZjaMvtPnuq92rCo
E59xuDx7ALQ/HmMbwYh0JCKc/yusYRGVWD1pv3q9dEv2fgpFCFRCkYRzV5dTsS6+a/aSkEJgcFWG
xUPvSwQimoeEOlYReIyXZYMNXidMaHw3lWEJ3u4O+QklRywsAd+t624CMyZLIbwfMftjaSq8B3E/
wesggLGegChuR0cS/7H7ItvKXplrSuUNSmnO5YgxnGUbbkQMv22VHJ0HiYe9b6xxyJs66qS2bWBc
dNyE4S5k5Sa6wxFLH9zo8Ac2WAjRxCNmlSZNL0oI4FikjS+Uwr6M9c9/j/StijDIINoO1DgYhLQT
CkuYJJhSPHJ4QSdtmZaVWb3XUXcEPDhAubndcGofdc2650f5swW7p5vD+a6hszbuTCTSxrEuuYTZ
t3Oiqsbs15dtYjuJBx14RBqIAmWUP3VC11h/1lP3zLWuuwyNcmYYzrK10/kmx2EOuLvFxupR4k2V
ayIiOTEw2gMp9YYBB5FhbpFdfwQi2dUKpAxgLlZOYZHBZBXv94Nl2gaQ/5ah4GwmA70NRf+iKunm
hiTcIwIIhId7ANZXEaX9uZA1xYg1WxzKVw3i3uBXNvyoYPLJNULqnmcik/btgBYlG7xfFxNzl0Ha
BUuSp3bKkJOWSWH2WgJurkhjqFAOxUlobKcqsnWcWS/78e/bMExaocHxggjZhFo83d7sXTubIhhY
pY+DjXGBt0Ubi5vfsUyYNwGlF7+x3z4BeOQsGmyy6Q7MggALICyMNHZDfcjHyxjCpJkBCfzOpE5J
5YTvkuEOHPc4pbZchwppyHGF8fDfXCEAcVL4PgWnrzRuZU+b7qzV1trN7TAvATflT8pQO6NOgA4J
jShWVzaU++ekgQ0IN8t0Ik2+DafszA1Gv5gsb5Bi5eYvEQeIiT2hkmx+xRrqNBt504AiRzWClc0W
saqvtOFk0r1L5Dhxk2w4/BbJMgWif9o4czBuQSTMldQZIyKB/53qv2DMLhWZbj+ofUPIuH7Xxq2P
Z/1XDwpUov1ztJSbBZwNyqRtciAGc8oF7OLx2p1OfGNAJCKsSSWCJJ2NvAMjGVJhMxmECiMxtZU0
XHrpY+T/na5YNspcCG2XsAvQQFWdzELW3l1L65qjaWPbZmJc3hzQtjVgQ08La0AwTb8Mq5VQuWYx
7GFwReQzsw8wBWLKl1hcTmwLaslszIezOXBg49Vko30YNMj5cuKRNhScZM9X+TMmIG9+ZTkOsu3o
zj6ZP6wKvZ6hAiJEkL3pCYCEYXfSC8B2CxdL53njk+wmjL0ApJ9NP0Aizwcwtwans9EF7uMG/o6A
cX8H168RiGKER+kgFnGLsw+xHsKFZQdWJ77YJbjO/9ggtAFrQ8KvjDeiKQH7I2rJ/e878YCTh5Qz
W9yMdzkzRwH3D/Aukp2PV/gCglXR+eJ6B+TUqsV4Gn1BphHjGHa07W4QY9eOMOBkDLV5vs2y6KZy
8ek9jcuMYMarNzTMDFBOIEti2W4oC0idaVXqHtZsrLqtVpeFOUpoICW2G8lgXCsr6+gpuOZBvwEU
FAhepMce/40vVm30lNVHNXesko97+jt0scOXPhmdsgun0XWRQwOOAc/4SuQLubb51daXQC1nt25w
Uo6oiBVeDF+saEnUIiNrmRWeWYNa4SBUx08o/K8GH7r/nJ3n8rVaWXg1rt22SRSR1RvX1b8hhJEO
Tj/C4eodlljfv+xuu2fx1LkIoqu5wzyJdLhDkg4lVcttM0ey10K7nUq0awpKmoCE7z4yh1HeGT4+
0J/uSKG3uNXjjKTceU/CAdfBACrNLUAJs+40FXvncDTO88HsoJ1O8QRulU7gKbnZX62/GJPtuKIj
ILiptwnSgQYSwO+RBdJMrKK/84BRTnRuRe0NPZa4tz/LaGDFQnsdUyMOUAGjd3ec8k2AyfOgbgG8
J3PYol93m41rELmsUV1GNTJPwfA/QJS+ow8EeAZv3dMcQC+yU0grH34ksW9Xj+1WOFTcKc/wltge
UevH9akoORZjMWzaIG69uPX/qrLJo8GqGoKWnwcox8rosxfRERk7q3sb2qnUKTLXFKWaVa4fwEz2
0+nJvsIIjjFgIlYbNyugutwARNwB9B9HY4QMnfAMNpW75QU9vYm3YKK910NS3jlykK/M9NDmAa7m
lRXcH59UwWLDVdZNQeu6pYCaZfazTeAfGP0sJpv6RUaxxvhUKlzw0OdRW9bDtVil8qsj82kFS4Vn
yl+w6S1ol6s4XLKyqpOvD0Az3IjWLy7nnG/fsl/EsRAEV0FL2SAqMP2pw9whOTgwVXePzZSZMnZH
v/8nfoLajamJlFs5mC40bynNhbGF2eVM5AIdczx83T0QbgsVrbX029PaEgR1MlPLRvBZbcc29iIb
A9hAJqjS7yiSZXTOlh8+ttNFhGogkABUhQETD+rVL6w20Zxsn0jfLo+Hw1fAPaIhqyfcdjkliWSd
+EdeDjUNEi9n4/T8/sxII3S/7zH06O2iBM80SJ9s90P3jpYxcH67rfiv+PKvb8No1Tb5DFX0aT10
jtXSr8sXHZ1zTpahayOq6OjPP0TUVEFpdHphjRAtXFIPcrM3d7+aik34zDileo2d9We/7egG8xib
VyARZjtK0u8vWNhWYJICGtzH6CRr7YI3jQ+DnwNaGs9gQccg+kI0w01/LDZCsoMQcVUr2m5Xx6gP
EHU+3/eiH1YKKnSk6fqsK6J3xPkH66X9ERHsc+FMxOeLtCXnjlAQ6lKwmnhpfDPFIeEc76mEjFxE
FXRPLLkNudAjSYoEpj+P+tYznnxXKGlBpHHhCvv9RLo3Eu4qgSaZLaB4+IsGmaAzneMpu/QB1eUu
5Nv8pAov3wR6MJH86S9uP281yq9ey90/ARvCRQrUeSqDHHH8ElQL4rPM1EDS1Q84yYv8rQvn2wM9
ABhSNi1/uhiWXOIjRwfVpk4i1r/fKzzhgql1mE1TDxZm2gtq6IcUR8N90zxbiVebOLHEAiDGWusV
+Scoherp6USzNdghG3ZyyN+xbLC4YcvPTQuZDavKwGhXqKwclmCm43ShlQHNrO+b2AYSC+8AJ7o2
pApbdhblR1SCV8RItzhGRZxqmVJhlxh1JnWSXLrOrnAKaUG2BoKzJvbXNnOrJb00XS+Bj0lVikPL
pKRj0kVHBrXmxaaBwKUQE2tXrGJAPg6/HflNDDsxBonjZ99Y1a90QUMsRAlvlQ41Vba1eBmUWCbo
UAPxbZYz7g7QGX8MsPsTx0s/eVKFSBauVOr6F9tfYSCotpwmZalIY0ltUoNvfEso6aXGFRZwcFi6
DYFLQJZA00XXHM75CEgSM+X9nzipEp16+lKP30ZkYY0znUDmmWc6PSVagIBHpaI2XM4S6u3LPNYx
39TcbdK9OVRLJbjsnLaCM1Rgb6csUcVwqaCw8swl+/Aojh4DYjaXabJQmafrLj14xOmhkYiFRlVr
uwr1KhTRi6QC5TO2JAm3+WvuOslhdlPWbBn1D4PqTvTcuQHsyYwQrBVxJU+t3seSTVFUgg4aZXox
3SUHRm9g7528ZoMD759IEboTv3dcoT6yCTSmb72UnX36YMJ4oEaOur/JLR7DT7CpDMoH28a1W8ij
S/Uj3bnNTRVVYm8x2q/jt0UVgjz6cDkPIMaFN4WDF4+hJJifD8NzKnzx+WheUhCaAwfTbl5FdtBq
oDgLi3bLe1O5ipPoM6DA2HqR6h0a0yqAXEgCsk+f/VSx6RqWJtdkeITfzlATiL9S9Y9qb8U4ON6z
6/efH84W7yrToeAoGr9F6yYhNzhKsobuFLRtU8aUR1Kk/EZZmZav2TaNyQE9ohSQJuA89mHIngsO
kW8DR7Fy9gBiM0IHVv01nhU7NT8srUW2zaG4b155mrp/kYvJ8R7R9QuNjI+A6zCXHwh5qCSfHQgV
SOydsiOSoUSSFZoy7eCbFEsQdQd8LSe0nNKpkwZviE7Fm+byFPPlUl7mTv5S0fCO4H93kXjFe1Ai
ztNKV0lL2trgYjFWoAKOuc/BX32SWXUOuHIVIxOv/fkdmQowgwCIo6Zig/M76X6GbSTvMxk/u8hO
Xq2cVC7yxpOa5H0Mx8Jbf11l0C7INhifmgrmVv+t52H3R2IwD/W9n3A9zSm1GUR72YHqJNnImHrZ
E2QtbkYuyeA5TEuyJeopIxxhC0x4Ujzp/PBZmcoVeNVqLSj2sgouCxfTqxAZej4uDD22KFtVxPdB
EinbB72S+oxsM9JYGhjomalxQsaCP+aQ9Q/rvmI7Q5nTGUzXh6wXmVVx+wgfdAAhCmdOZfDjBm6E
QPrXtu7zbIvTkPh1qFbIt5TGcOKiFsyCUzhyOGHI4kq0tOiTpGBeKAhfT8ktwJUvhp+BrXqxR9VJ
NyQUiG81iEetYhXgmEhVd5SRZYBDseHr79BR1GNrjIBiCXIvY2JEAlOX3I+rAwN8Ii91ZqU0tOsr
K4WUi8GJPpM9llLNNqH7DfZx6ruLOvumAA5UZIaKAhO8nIP1hxp81DkixNJ7EKp7UZqPPVxlHstT
gsbRjGyt5fFW2TfAXXkb48yX5ZLoMBFvwANYXpIWy7Rs1RSYcVUocjg7a1TuQ3JQ/EJAH1P+MgJR
CN6bzcPJDJDGgeNEnnsgi7894tI19QGkx+E02k1O4TJYNQKyQctBnK+0CTopRrysW5+aX9O9m4tT
eONszKpqReISwhiw3HJ/ifCmryC+1rQkcP0r5qLyOFRg6IEm5p59o26tNdFeHpStUHLSqLZetyvA
3Ph48hvpbzZa2R7aB0h/BTuaALkBwEfx/1iyUWqMI0OJ2D9ZcMkyd3fOpBaKvQK5AbdD+i48zM+E
+Sb91w2r65r1iaFTBuHUrQQ8XQFNLBJ5Ejbp3xddP3iA2dCypDV8pRDjC2/iN08DDEijOB+0wxaw
kR95kL8hI22p2Z6CC1RirbusrkN1Tl2K+4RtEiUbbOlH3X6hfpIn15N43mbAMf+XWzGU1Y7JMRsh
583BsYPijPfcaevzUnXUU3MM5RnNMzxi9hHO3jxcAzZsmvZ1lzNv/hNJF3Z/ZRsxs1oVs3PdRXbj
MnuXbfNsWj62WHPMqE+ZHC27J4CYiI+K3SXQsOgfNNnkogxWgvDY+x4qLqfzKbUtFqGCWu7FBtVd
wfu7cF7s6rYbgB1k3PipNL5U6iYAYDFVmx44dgjGGjpZCg8YRpqPtbJj8EdsMW1ITBnM+mTyidHe
eDoNKJBxrbJuAMJlmHfHAahbbMakB2nGBCgDCTrvT/DFHayczmjSyuHnbIaDbBQVJAM/uP3y3Sev
tXZKm+CpzldbTCVf+04T8p6ky7L+yBxpTcO8ZaosQN3vBru3aAAp1IMpARxAf60j0hBrlmCB5s9D
0YSNjGVsIJpQULMYgiurNDJQKn1i3tS5fFVx55NoC9sJcJXKaiGj7qrVKVooXKrcswrcdeVMZgE3
ypdUSuabT9C58onbAbGezLcuBRbynHUisuFTsLlf1rU9gitafP0kLGUB+qtrdSGbcGpTeQ2jCG89
KON54De1Olp5YCng2A4Z0oQxb/GxNX+UVxT44V9CLjcFHUrQBQW1NuQGJWuNPi7VLp6pmv1qQwoG
IdT6lF4wZq9tJMC80lQMvREy1rkC1SA+HpeszSUOIfnaHTc09lU/19vxhIhPFMS86YV1z2hgKsJX
j3oYWSMON/IqZowpL6dZoA6QVvdPjVh4iVVmDNmDzp2NwhpzRBrPi/wP5qvsVqWj8AGi5xtjuLSM
qO8NGQe+i23c7VFUmnmoIQ/Z2p2J56fTOGGUDA8g3agJXR3Bgiwkb0tFNcVCMufN+VEX2DwpFrQw
Grt1ooqZ4eqNdpNBUlf3tp7Fwkm9B0j9q6/FfC0H+7M1ls4prWKS/bokKPsdWsHdFLD0Uv78qhFn
CYOgP/l+CLYlHmA+bOprZYh19Rzk/2cd0neptzIuNv4Z8CMFa0EmEurltrC3See/PkKtwxdaTV8r
pNaETJCw3FW8eW2qQ5MDHf9/3EY2tsL4oOTho3wG24/KAdYwc4jdYAKGTIB0OZxLrpPNySj3TVa3
keVmnxcRHyXKPvkVmoZU+u09IjeQcbU2oIK9ibuaq6cOvzmamsdrr3aKWrg+ozD4S51uV1M/3m7X
LRhOc82sHqoyslFr6kY5LrFwo3Ouie8BZvKXmxR4TdoqXV73Tag62e6Ngf/Qh95EilLTlrs2tTOE
lsloS3rIjVEwTOdrBEJFpSnqqoBbYnUQ5x3RaWfP2vPWibxG76FQt2vYnlKQDfKaSVmc25pAxxFT
h+wictuqUbh6kyNh9dfEKAxGO3KNaXZ1kE2CSyWtMeWLI7KqOYEtxqDPttwTJlaVc8Imr+aLxf4P
U8ZunQnYVxKpXqKAHH6QxXHTAvgE/PAeqZg9VS8UosyUCXWOrqx6w0n9HcI4KixeqS3VO+hGloUy
CZ7Fbf3xyLak0XxOG/tOAuMuxxjMtUgYfZnz0UibGY3/Kik2wYX75ogDWHyQTVu9Jr9093H84PGE
BlFm+A2K7DLtCCCwlpRCtvV4eTU1443Zud0yQRKnGf82MW74wh0124Bh13Oc71FOD6F9eluXYDzj
psrDDrnuW+2GuUn3Wmft6TnkL9QjqSvycPmdtFgZsMATPSmG8oZx1RYZVPNkogjJ3Vk3S54T92/S
1NjsoDo2CQlrqbhfuBMMT/CQIJ1B8izUfoQQXdsmwf9pmQIW+Fzc6RNW65yLi3GZ21pYjhZa/B69
0I9CjpDH5CuUR2Eg2ld7j+TIZ9JNRTJfM+W4ODWQVrjtJO/TnQpgEq/aBPdijkgPLb4DQu0xW7xK
YzEZoGGvR2zUeyU9hlGd0dMBQ5cWCo0paqgSfC9ZXtVf8RPz+AnZDyzP5RQq/OuH+3JMmYvLCQXx
4MauzAMrY27EtqBO+Uy2Z+qaz4o3Rmlg3SuYB+crVc/Z6h/z55GGoUMYbs6XmSJjtUK8NoPKgZdx
sfoDfGGQzk8HBZqTsuCyrvkgShElix4L7p709s8QsZ9Utw5osJ6KDmtvVohX+lPARBk2fYjDQD3j
AvYgMX/gyKh0h/CjQjc0H1B+JP5b3f5IqUiAK3dPGFpJSew47XGLpPC3EwVkEXUu0nw/0+Rh3XXc
ugN2b26nNM6opFa9ml2HQ87fVVWymx9pwH7M00dMAhWdglcEBv2qHhPVOIdifnfUfEj4Il6YjNXJ
uc4DNDvUwWCBfoyZDYigfCeDCPD7XYeIU2yrsg2QHqWsbbnTlVBApVRcsr9K/NbhnjVIImsPTtkB
62EsUiC1FPncf3qqSRDn1MayqeJT+2c4TTtCnMFz3ZyjB0vHPiyLt8FOSc4Zsi44JjnTiJ4UscLN
pEf+/u9AXTA+5EMsRISeAudVSYk6Ss2KN2fKsvCaQnj+Ttys1kVRjK1IjEhVij18IkfNki1EYEJN
l/GT1m4zAt++O9io9v2Yj/6MmWUCHjKn6c3N6AO6I8ShQbpjgIupdJbOzcf8gmWGpcBGY7HJTYox
tEJAzdyGpkP/pni+RE3qcjCEUELdTdXc5ZeewSXIq3iAiUJATys8cobkqG4HvQrI/FpWyR+oi70N
1PKf8CtdJolD99bMCkJKkXWO+/HDnAKyMij0iDuDPUsHI43ly1P9AA9WctQe5FRMRQ9/AMuujYiK
fwYiNlz9Oiv66htfjx7MA2M98MeQdXPzl2vFU7zRDpBIVigoVEOmwX1z2T98JIPPwI0m4pKtfsLd
UwedWCBJDWiw3gC7iiFf0Zip/H6M6PNb12HRE+ZVRpsJFOuuF0hjO7MTmufkdFkM6xseeEzsaPzK
ftHCzQsdx2DZUuIbgfLa6JsTPikYmVbHyiOrGtlxyZXVJNBJPcvA3k8mhjeKsETpbsUkXZZgUKXK
xU8xRJ8+ZW6o1GNQBiEAcOvfmfcCcHkEoQFjT39vIMnmcFb0e+nqQeewwakNy+/RMdAZsJwtz5gg
ppTyuGwsz56gxjOCoJcLwzbgzrcmmu/oAg5wt2hffK2F4OyrafJi+zyW/HXXf0+dtrpsa3u5uTos
8zEdk6Q1IVpVN0HELJ0HSqbWTq2aqqXNgbQygOHSv9btyimHwBtyQq9VjQi5FaFvydRhRAtlQ85v
dr7q6N+rJRSi7zf0fnzYBr8sAo4Go8fqZv6zsZp+bbSEI8WcmsAhibrWRJS4HGpOrV5fK+UeYb7R
OBF3u3rhX47ZfoRL7F6ZVrVggVJfqMWQw+Kw/A93II7FGGGZigAidsFV0gxh772bZeb/M7+rJG5Z
KLNqG99UFIhZjQJeBryzHlfZUOTfSJgxUqtExfTb7GC3wHmzirhIc5qlmCF0k8AV/4TAreLwKOkJ
sLfphyi3cKsOBUaflBMNAZYkLx2JCn+0zUyrjHv5DhzpGKl7+fKvL8xebbOB5eMRc3gFQjjxRs5B
td93Icf31MWvndFYWNQHjbU6wD0EeazHhGTyxcZ2WRYL2CI5ZA7asK6knfNUXWFZjd9XYnu2pZ0h
20vDEygRCCrRau71KRCDc1BdBDT4dql/U1HPHGs9O9tiNkH7RC2t+KzulHhuVCCRH4dwoF7Mzefn
+mNEst8GYCI8Uwt98ihxKswtCfKfMVjSHawTafyhaccfSP4nojocMLjw93xizd1DMqFxPpi34GWF
ARJ91ynWzy8rcWaSWs46aYsnIZGIx2rCkNbr3wocLvTA38fKzaYBGNVo0A24upq3pzOgrbt7sJB/
yzVgbi9IOTQqeTbnm/0+pEYWHKSxLUTp0PhmySgmhmDz251vdKKqkCb5uMq2SJ3ci2Mm2BUTptVi
/BT3GxOOYnfs/jAaN0rJhQO347UvWZaArF13XQQ81VP9XU6nTPp1czeAGu/m46zG9afQwNgakW3Y
fYUXByA4nSMf7/CIuYMnKYZbpTv5lMVKa69JspB+YKKUa2X+J905uMLHS/gWA+b2R27ElmPvKtN2
yJtQ56mGs3gIB10LhEvgBft8hMWu7iwZn8w/FdeZk7nUyXH7If6GxabdVeQ4Gbbs2Y72GgcSX3cT
ycMLDdvZrmmny8syww/eXNo5NTWNCuyQhMs8B1Q1Zr7p191vLQliWKmSBni1sloIkGruVEfAW2bA
1UjYyFoo5lXn3Y5+bfHQ+EtKvuCexmca/JX4264wyFs6DAQryD2t4mTKmvbdsOkh+RcmLZPX1DhZ
rwgsxvrtHmWHzsEtyEkAFPcLoFEi84Dkir06BuIU2FrhWppJ4w+JmlIk7dAlXOK6bVln9uz4qrAf
gaAlLWTKQ95AcfQ3zb3IZkpK64AV4RWkrm0LaIWe2bWlrBu9qp3VEnojCsdzmqfN4MXpbgVyez/k
psANxhnAO0YxUbJtGeGLcfEvXqi7kXDYhcdj2BXQ1QDQVwQTc4A2xX8OGTejFzJUcx/2hQKybXVv
lPHSfDyk14sqKF26Vl/pfKeADtpFZk3xXfF7kZdhE1/VZ7eAsJXs/kzxXcoDnLN5BkBcHfv6O6rF
0x32wH/jNfk8N4TAfvBIsl7vKK2bETLACr+2y63u9lpjqa0qzKj+mcCymBNFShWvaxBvbBueuU72
Z0E8YxFUqQ0YqYke8ncBjZPMzR0yJcRfdG7c6i2mGJE58PXu+Awc9uz6FIbezoivmYIPmZPkRWum
btSLiJkjOp9kBAUFpjTxQNOcKNlVwklnjzapkP97xPQZtOPMrjvsQ+9vVihgjZu8EpxF3kG9EkLR
MBNk/UEKmUtl/F0hhYfd4MVOU8LMBBMFj8rQRi10WD7TMnb/huwPQ4RrTNpOsuSpbrjOz3yktedu
T8kqrnSq835LFjZuPeJ3CU9tzjspswvi+j/pafBjSzvOPJt3AmfpBd6X+nxch6jv+fSsiyMuwKuf
NbjpGkl71mMvTDyLTfGfgei4S42oLL6Bpp56y3ON0OMejF0VxASbM47FxY0bGEu2iugu9HJSPaSq
J2fhxEpgp1hiSIt8WCdjoAniudTdHCEYPM2teE4tsmHR/e3plnUNiqJUY5aT50lZMVMRGMx7nkZf
b9CQUazWgBXOEOyxFLuaSzJoZMfxKpjnueTBTGlmEuf5fyl92/EpSsifHBMlUE4ltDywMjiitv2D
bjrZJXV5daEsSDmxZ0RjUfH7jXmZNPggTnJqGvACwF/bq0A9gfTL0rjeVpFx594KMwzfLF+gjiKs
u/XjlvA5isFzPF52yzOuFTiXNpbIIfnBcvZCDeEusR/SFqF39pFgT8gQWUP3S+22Iq6UA1Og0GEk
ie7IjT3TOdIhA84GNz3Pp1pNxdxUA0aK5UC6W/YEjoBgCFP6MhTSGeAmz3foZstGGQVrW4onpUaf
v7QKS+zVLlIZQaeKp06OAfX2lMNQ18BLzNRAnfPlVUrJyfIB/spjzEFbWCrgNJh7ZBc2X+1B3jED
e4JZNc/i8kCwEW7b+0EspDY7e36QOPZYkhsWyKTkdKlr4T5ByeRmW/wzIupAz60vQg90T0SWG8iq
1d5ntK4ONiEkFFfMMSN+pDwk6rcXeFxB3EdlIli2iEK0IAwXLWDo+os2ecoiLB1dpKuQxCvq/tmM
GCKS1lKOQyTof7m7nRKclTkt/g73AR8pUdO6Fqb62LDXMbxdAB25VVatWh/e2VvffDEbEF2QeROf
w6U9TOBs/pLa3iQx2XR0PI3Ex0DmZRAv3EH56BzuesaOKEXoKnaXtqMXq9Ksb4TV4IQdZAQei4Qz
ieRXml8sVybXGhegEwdRQzhEbYNDT3gY8ZXtXABYZgeq+Hwfk0uQyxLbsBNo8maxSz31/uaKaf73
j4CsQiBk1pBIz4KTvjkF7SVjiwDFcoay/TGvGtkClos8iVYKkj6iZmoCzbsChasDAoN1olJq5xcA
u1cgkCcY4mHQhQkwB6nDxW6rIAbUXc124Z/ibmIEXn3XoQAK2JvmjU6PUhi3fKJKPP6pMLBKzK5d
wwfOKUnobfescIne3MfL4m/axVTjA2xcRYCNp3oiYf1CNyx1Eq17TLXiJ4/YqeDVAOaH8jW2jqfW
wRM6lvvgCoUgdobjX14ao0MLYcCmXh5Ymclc6Bseau7jdW6YOqit/YIbQ5B4ln3DNIxjff5gsn9q
auOtXavYAyQhOhvqoDhis0cK3Iy+o0Wz20IrPd5gXgXPT12V8XTU4BB1OFC2mOkknBVu3xXSZsME
lmj/52d4Yj3EYbqQfN33PYZCNK7PP1bY8kiDZU8ap7mZSq6uO2OD7YDgdid2s5rzbrtuIms1tPun
QfigBizI9umToles6E0GgGpiR5QQyCnAhCEbfzcjqNjt3M2mKuIDy6qy3KsTiYM6XrtASiV6Y0p6
NViAdurW+5vAKcqnrALm/slHpefHvhKKn7Z1pC/yfDaPjOtm+GyEiIl84HPs76BAt3139XPPn2UX
4CR3nLjh+504JdkoaOnYJd5k8zLTRr0FTqM+nPNTJdmMcRZ6x+VvaMbwemnWCB7a3EPQe7n6+8m4
JLomKQzSSA+sQ/164h9sDCsCdcvneCfGhfF89/ZyAlj4RUOnZZy750oOL3Q6Rza4x2eV9ZxIxU1o
LqClBC+lRsfBv8vsam1d94YFmHTIccH+IdYmndpmgQ6DE6g4g4A83A2EXxnnCF4IaQFWFIQ9UUHs
Vdx6qeCaMzCQLWqdHZRltYNYeAxQoviYqyldekTLgff2B2L8YcOWRAVspUqzOyUUupMADkkS5NGK
D2U6v77WIH8errd+wikurLEvATx7Q3cOLe12yg15oCQ1rX1DIU7swMdt1yuHLGEP0iSVLJAFfvWt
nki/BNRMtkvMHviycXQN/57Ch+0xeYwp4HglwrsfIskxmuQfiXMQL2CNxMkNU+Ht7w4s1qvLjwPN
DltOMnckEwhxyA2IEQX9IdWIHRuPUlNabz0YDhH6dlxJNy5pgQ9r2Cv/t8rj0tAmX7LN6P8vJ2yB
z7s9/TIHEyFR+8GqOZuOiC11gmonftVh1KEuaGe3xu2OUMTYrxrBu7AaU8PTNCgv3czq2M5KBbLh
AkG2BucwDyPJ+12WGWUN4krd8dWlBkGHyTudVkTo1cQSdEzd1bbE78Fsap3adN3BWjdDjK6hKQzL
KqMkurL369Ms4fDrJTp0bGd9UziVAkE9ic3ovC6G8HQj3YtZjFDv2KD0YKIaeZOx3VxjoF4JVv9U
Uz7ihyMTofjCD/UTOhSVihhoKvkqNCFU0Cnr5URlmCpRb8NynxdcnNHe4gnlj3agINe7ywAZGoVv
MDswKNUzlP/MFSv9blwxta2JqqxLpa37dTdHakTpQRm/xAoG9GodkzJuDEbQ1ubwXsdiPFusogX4
pzBrrNj2NpHKEU5mrvxBOT+NT5qkRSsA0gl3som3K77h+ibSH7sL9f/XTRywL0NzIHv47W0BIJpG
ANbzlXDlnhZWweCTTeWl9kYvy4d8pM3HXua3hhWgKRitt1beYfmui/pWYvCVHImm9wHEVFO12/4m
pgeQMyL/PxSlOO70WRCOJ60zThUxutyehTyQsATQWkWcy/dzsdAUzcHAo6/bvqM0ZDVXnNb60wH6
v8bteHPfCebr+hUUYkPH+hDTlfSktdF7lS79C1rEZxIIZ0/M+MXyn5dQpe8QvkplO8tSFa5htbn/
AGIEuKOURiq8SsXxYumh9KXfmz31Z73BnrjvJ3G4XzijQIxNSulZl7c91h114yZS2nnL2+qS9Ja9
Nm3Gf57oLUwreDXmvatl9iJJ5n+bKDPPZgrokBHiDorbsUcHair5ad2GSCNXGg0H66XuXIevqLAK
LEJMBhXDsZosuBYhpn1hsH8t2x9+KLMFABz/ss5yoFfB5HHjGle5B7YVxiQlT9kQekBxNDD+2PxX
oLLQwyriIgdgzSWoQpmWTxsNAxKTZeblC7+vrIgtExMn/4dpnPYe8jaDANnYMCV2IwWkOdCeZTQ7
PV/zUVDdM2PZzn5jbPuowm+5ZTQSOQmKIASxph+paeYkxDJl6mkZ7lgoFEZV1UlVn9duSOXL1HqE
AnACKnTqZi6r0OzZJn8fdbQx/LOUzkgMUY4/ECLYZx0QpP00D55HSYFMGzWQwC45OpXjJMPfGL97
/IR67VlkFIeDX+vnvAo5uqQeDG+7bMdgAJL409Aw9A2ygbhiVqs5YIrlE3QIo1WY9nFngegna1/o
D+3SJ7KKXRO5SIlYMM64Ze/TXtxAa1GHENGlvVOYZkEuaQGRqoUJ7spEorE/Om4M91x0G3BcpcyH
BzF2wb6Tjrw2haZ30qOV1AgF9x4godnqkjxOxzBwogU1LkbJsX24eppwgZe3+6+yF+ztc25mGIVo
A4YZ5Z9HOA1o9oKAYu3nTBfpKu/T4iwjwHAfyCmjSkmStLpZ1hMzt1+SQzgT3YwhxJP7gpoUBslO
dB/3jawS2typQFEFq08QNHsvovMF/oSvcU2l+/VkZw6fSSMeK2l4ThWxtUk58R8oBDN1xtUy3OZ2
i8+eXgB5u5cW5BrijdRkswIfIsVjAxEqLEHeBmpaURubRcv9bB5lR9YwcwqMjfTzkbrO9PtD96Id
i1FPaNMS1ilVs7esQ5OV9iPnCW/FX3cxQGieRoxW8AZlzaoG2pI0HJzblKtq9EIZkcsMnoB235tO
3F3B+y46R73TRTopdpwHvVetZuGZQKkuQfhzE/kPsysY5U6oJZ8aiYN3jJIJ5wTOr826fYKF6kT9
kxrPJOQEpJx80gKmCAX/xVL35WG5W2al0cMKW7jPXAH0hP2PRpant3LTa7sXJs2wbNdhW2a9IkLB
kgUYsJ096HRVhm9tcFvTCod2FpG2jeehGukQI6aK536dzo2METGcPHi8G2fjXz2quIU5EyzCshxu
YKOOD0EW891lmsfZCGw0yHl1RJc57wA0FYhQOApaclTpFof+RDmADD9rpeLFV3y05rnCfgLQg5Lx
yQ0J4nPF0RmorGrBJ6uo0fGiJ0Xj6Un0gHecCG0A4jG9W6NFpcEVAf7shgULcnmOoAHNwNq/bk9I
WaJlFYCooMW70Sbyrf/rNJI5KEu9oOyBTkazreOMK49YulFFJxii5uhwcZvnZE9pgKgVEk3hFByN
kJzsWifBdTYFg8S/0Jfcumu7O1xQUcGhRqud2aWGhYmKevla6lPQo4EquNEuRm30dVle/oNBYxWn
7XSSuFYZ2BkyZZ2tF6G3WBuanZLuEBP4nWhzcW4BUJWk+C+CVb8OLahFFrZlXS2x7yF3WiwtON+8
4eeNSg4F39y7YvLqYUOVEXzlV0hIDAWBR47ywHwb51xKjfHvwP6U84LsAKMVgwwW9Xm6+oxkR7mT
+WRmNzapM2U/BtEQ0Aw1WUOO1vtNeMolaYcr3Cn3LFJo/b4jPPThI3hqjtmNEIOjdY4gl9jxMd0L
Sb7R4n0NfxCd1O6fMprDqUzpuZcc4rfiB+LtOTYF3kvwSzrbdVlIabnXQWoQQTSEbrfAFNpuovXR
W/ewfKyj47rXL5TiO8L292SKUaEZp7OtVixMIhlqq9LgNzjRcE2ZfGQKs5LjEhUpPaLjOzFlw+hE
x03Srqe5g3H3rv0kyCLKNf8gy3HJuFPCqteuTxn2N85uhIGwR1k3VaM7XhtBiDTRBqsUumsczY+S
v9++iAEE7TJNFJhdK087aK+aNKJK0lTipgpWEsUe4dzHE73498UMkQ2cUzAa1xSks7Mess0OlHy9
BkgoITz+pnuiPVIuIQr4KoOk6R2cANnhmOASpjGVHMb5J8kzSY5dzKxoJjC9uzKG8TnOv7f/Qthp
fE6cjdTtKohrn1i/ywXrpOLcSJtk1C1ouUgM091RKxVSs+G0iXAhQjs+M0LJTeiN42MmNFCFpnz0
goQLxs9x0xYdFaCsehEvvMC0tgGjJXrcqPxNLIb2kVrjFE0rzuT2PuurGalmxL9FwpF8kUPileqV
+CQwIELrYhftDGct1HoZI6M6Umj5P9Z6IhwAzvLzZenXE2wYoBwag8WZOSAM19w8/DYn9Mr5XcUi
5fcvSslMixdogKAKVjyEirrXVjvjAwJc29n2i9m4jOJG5zQ+mm0M/kVgftPsP9ISllbN3i62YvCb
GLxfU1gpvsv+QUo9Zi0/8HFtWc+ljWRQrEQv9pB0zb+moERM5ct/e/1lRobe2npTRbPAbuc9lTcQ
g6/XJnuidRzgLEcLfqioOnL7i4RtLJuKWpOdiidBNEQ3SWgu5vv5y5+TmDrOvXSp3DQyD8oVa94U
L4KkClmnbBZgnZdNY7D20BooFjTS5yHWS61c+BSnpLt0M02QxiqDCRI87JZLAwlxtKWovgemBSv9
6mDH5AvWGB/LdMoe38I/vFq8xYfOVf4227YVNRrAzLjXAa8+UOx4J9qYgvTQhR8EhHi4RmN1KKTc
nLZK8pStY85GMMqw7tGjDjwlQaNpZ1y4ZOl2+cmqVT+15SawW4EkQNbavTPSSJ4ucyyzPxoHkVP7
ihq13tJWdSFzd9T79gSB4gTi/bB+j/ur0Q+49M4/QEkvl6TF34GOPBN4EysY6zBlcASEYIOQ0UXN
NQHIgDa+bYKSG2UYGuU6X+p/Yj46wKmfgmwtxzdKdMQX6I055HJ+LGaFEAhS6xpPCACsCSini0FD
8V9evN6+4+eF7oH/ct0VYyllLE0etDha1g6Aw71lDInPh/9U5ZbjCGPjXRzMulOuR5eimf/Oi6St
I/KZ5IhlDi3oS5z1MpwqaJIRoQNsAU5p6twrhJoOe6Ugwd9JtSOCoBbVe2qcWjZCY3OeRCQCdOhP
i9kNZ+7eOhuU76yWIXyei+eg1fFd2bRbJaiC4KIrTOsVfvBuBLFtdQcEwYj5i+w+2TfDwgr3PbPE
2zcFGIWNfCTMCkyt+FLlsKYMKm3jfyrT45nKGYlpCRkjh8L6pgTLwQWNA/IMNMJLkPhz4arwKuED
XbWCgKl275HupsD4sxaqIxYx4n2N9w5KGEBcG9Fujy2RH54AQ5Dtda3Y4uShrKGpqcMcq0e+mIw/
RK1dF5A/rjvNJeaKw7fCsVWvIb1S69gzpa6shL5rsceu6eop6OiL526AU2w53GeMYFJgLS+Ns6Ry
cVUXIV248Ws4fQcPPQSqsVShhzeqU7M9lpCdYn0WtLDElkObVyIssW8x+7xurd3/ut3BH8m/GLq/
mnFRhc7xE5xIBVcvKrHPeyA97E0iFRkIsQx/rE3AgU1bDcIaLPdAVHk++GLv7qfLIE8sbKGRZnNV
4xtp+7l0ZnAGQSZMGU3zSPl8MRhn666QPu9icC/uOGvKX8HkdPjF8LQb1PJ16L/ldXFOz4fOhlIg
5gbwIMJPXKUWHeGl87eW1lJnzkyxVAHnRHS+ixmtBrNsK9dR1sPPUx18EY8Ex36KjjF3zYpQJtxr
Nywz7+1sZe4n/rxUvmXTLk2QVUJI+aJFyROk9zMJJZ08KRRtIigRyi+s1gJ5e3/2l7WXux/PoSvo
kws8hwmsL7z2EisiDdEdaoj8jheIGQEIdl83Wg64fQLWGXM6oicJDBfrX+ntEildO77e5ZPe6sHZ
TjPlJJJxQwDEYDpMafJUeUS0pp0QD+dc2+e9flZHJ3DJNhtuvUxBzVgEb19PlnRlVSjwHyYcVQ/C
wW8Ac2K7qiqZCDHijZaV3e6rnaotJZ4+JO1f3ykHej/I2rtMeW8G9XdrtXo2YB5vVyx487PfodSM
HLVNxzJf30AOSQVL+TkytBY63nu1IdnVmR8SVir0irapiPdqAddQsxhUFbqO6scYXdXeobVD8UPL
ZSfdh8r7KCWkbSzlgTKrPzE0wWQeiYEd3qrpZxmw+rexLiolyL2JxgsySyhq9cE6Mw73w0IU7DRS
2FRvhtTf9UyVszAQt1haEH/LmYUEB1Ayp5AXWg+WSQNPZPlwa0Zf5nmGZO5s4aj+DgfnXQ5wHPIp
vj0gwaRA6QpMIqH4gmhFeTIWeBDX6JGHRVqpHVFC+axZp0C1X63QXJuFO3KLYdDSXByQpyuBju2o
XK7502pQYHtYAiwB9gcc2i/Dyk8YJuRWLZXCpD6gsgpX2ECJkxncmM/Ac3QZ4Eq2UPl15qNWHC1M
qdqPr+XY4CHzNUaq1PegicO52q/J66U0woV+4Rl5owPx6aRK4lKHtE9lgWkYen0+jKjSQQGD2qAY
dRhYkmuxlYTaUP4zUfndkkjSg/eiikNVu72vvsR7Mec8UUndZ0ZxCOJ9ZwHL8OrZxks0IZ6Vn/9v
6AzCHXmtk1u9X9bWhCRjfQ42pIMoJcbKObRrRuoQw7bMaIV4YlYUmTJMIn6d6Ve7pxr/Wj99sYMT
TmbPNkOWEiYJDP4EN/2FjmR1eB19BlkgSxutBRDnFEjzrYuNl3R2q/EALkXYh9meh7Uq4TzRRO81
gORATHS/rJdpub0+m7YD6nDbW06vimF+5+gd4CpeWqrNjGKuC3zHSqOBfIKDwFUQxY5ZHUzhR4X7
Pl36Y/B6vRIftx5WPui7CMhNquXl/DOt5ZSjpo4xWr+tFEC3jT4ZwNdwdZ/NoWqdoQj6yaFvNwoW
escfeKiba/wUFdEM9L8nEE4MyOpYsslDGePGJ2/vgoQAL9Ro87+ejzqNHyZvtMsCGof9xnAOHYHj
JDQn6ZKY+U1b9SbquCmqt8dI6O8HLlDrc6eBJam3guXcIFU7/ugENJN3/YOgt5TVgzxAHPxTkTrP
JZfWGrmX9zBF4A0Y9YP9qUYATOpKLHAoDSIJXqb+b4CucsmcrqR4lIvLJFzIUvgIelJ1s2m8NpF/
2QrMs/AQfYC42OrNA2/onvFty25PcELmJg+wt/XzOtPjzYX2anI3FB4869Nxcz0wWu8sBOwPTpOo
ly+O9rHquiI7Cy0VQ3zLqQv8M+vcq147ae7NefhjDiILfdHM2MwAgKsbj26U8rfXmkGrAxoWP5xt
2+B7urGyD04mHRv9WHZvFG3jN0fLfJSR84McqUCiSpm3iQjYjCGI/sWf8fIeXonhplIsjo+JFIdB
ZqcBQtyVOLjFodfYmV4ZfeEStwJp6UUC+TetN6jM3JQ1RLfmxqCp6OC1qEgV//OqIVrl9AovNapN
l76tmYBGqBq17qvMFNLwquEXXdMIGrDTXHFnWcE5iFbdaG6XC3iPtrRFoRxprMY99EhSRroCxbfw
VHHVWUU33Z2u6/L1HM9qjThULpeprOm8zR9frXDpumrjExytmPoNBdajMgxXC7Hi2SXOAInk1gcj
Swz+YVyE2HKLMrsre4zI3OuYx9rSRCQyfdJSjtoNeuhgoZeyTH+C10BICavIwMeV9vq0y5LEPFjz
8zqrzwsA84Xp0yTDAoGiCGlF25CkycCND3449oLl8VIP0nERhgA8mwVlXbKXP3UVFyY2Ck3kA1wT
d1MQdESPdAfCAhVNvdc7ts2xbQkIX8+ltqgFtuSp5Yxgkon0vlQaI12hshhzWuPjoYmeNCHyJBwV
P1VXpPyP0a6P+t01UETEDiQ4gzqZqlV68ejkWXUR0ddxMZq+ZsHHbhD0mGF2dsej3XYkmfiDk2Uk
KLjBRXs5kjlS5vA3qR4GBigOYPF3HYl48h/ZS405h67vazk4fBA5z1ruTpckdtLy//7uAf2HxkJc
94hvkXt41TFtYCtb97Q9BQz1lvCYhhr4+jjUQZNoDrrb1/e0pLYCJMgS90RLgJBWhWDr2soC/Z+s
FmfT/qaVzNACKDZhMZPZ6fZqe0EkqKIsPiIctsrMY91RqkAe8moBMYArhiV9Y0iJGZM8hh5Is3eE
y9Qw4mk0WDL+t54tYOfys4TOiiiDaK+01Lhak9QTGROZBUR2Pz8IBdNUE3f9yzleMoGEV/de3zbT
J/FaCF2vjiiblTYZytIF7MFyvavr0GfxHpbwLoyh49RSSINvmnBHZi5CT33sSMuf/VKeKcOkm8ey
2oqw/DGOauyenVIkVf6DkxnUde3mNT8hsLd6F6p3TLOEhzRm6GLDwmVpPya5cyMeknnakD4wKMZn
X7oedN7Ome0ZupbzhmCcEIxTNkKoI2qPKWiH6JLTfY1CFPSf2sQ7d8wyxk6MPffMUk26C7gpxyoT
EEkuwswizYyr09sUYbQfP9rQixpUghuUdsj89RwQ4H18iIa/qQU5y4sTj31ZT0EyVqkp4++VSeZi
/T7XpltFEWQOmtTN8hFd/Sif+KCk6RF9iSm93RwatCRKYeKkymeuEKX30CFOFMFva7SA5Y6ZSm8w
bnCSEBlgs8Rfu8sOmVMEBjI13qLdRTCr6HtYj9rSHejSdrhicMSGQe5fB5RgVH5hatPHLhkEnDF1
S/ZsFsw+Qg3DHqFjl9ifOXCSBk07jO0AFa2gBrA3dKfiu3CEnd2Gyxl5nCKoSicmwC5IuayWOqBT
I7zNoGDWi7sBF6KuENYiP6g2bYrjJgoDFHrmhP4S5FJ7JTpsdLkmmCqqF5/Jv3P+DTlEoq1DbO2r
pgTKvQcEnr0Wypn9zNmM5PsvSpnakUbTwYuC7WkAxkNgLMpbKD0P89xlrvw+EEDWbIBfB7ChwIZj
Brw3NGUtsp4wCVBxbUdm+HTESjVWIH7Yh82jmDGRK65DrQ/Y7ei/jsptA00ij8uBm7SacBk7Zfkx
I0+clv6TCopRpmld62Sp6oZRpdQmhzNA830UKBmXgwGES2LsDXgfLFEZRedlMHQkBIa85ERLgHYL
fqAT9SrEKLiCSSLqv/KqCf8TDF28RKOxBxdXbBHO5eKG9dbAijVBqWkglBK+E/NLfUfoeT+IONgC
e+1nn5X5BLmASOYkEIQIamnmfxQ43EW4dSmmBjxJiwqhNPQHxVta3luF+0EzUwQVbvd3bWYOrH30
nAV0J3YMpK554qB4K7lueHZmLKBkFfkoR9zies96wfc3TV17fDKZWtBNiQB5OPwlUl47qB69mpUQ
ruegbBK1YEwOO6pVQ1Eu0jsGGtZgcDZmfr4IWqMXyOyKKNLgbfcKk/z8xzNMdWXr6zbmD7Loygoz
qjRmYCk/EgGfZFu7CtDHQxn+noxA2M3tBikMQQogdr6E6kLX9YfDLyz/fZfoWeRhefC59YmCuddD
ONOsfiUcO2BMQwVu8SUDmgwuNBZMS6fSbf44v3lZoC9og6XAVuWJIsbFEQYsDcEJeJaSPKynVeLi
DNzGh99DDGUMI736MXE3acM8kwgVH0vfHqMB+llN2zXIgpWl9YLM3CZvhuKFD/gsVGihNR0iwQiY
PiiO/N6LFDE+l/VM3/3zm6XS/ehMp+KnHQSg92eX7p81l3x7lDNcHUzUyLfgWrnQn5X23O6H2FjR
vgNA732A9+1FcaWhEhp7rk9J+n9W0f2kvPBKE14wHs9SmheHqiHqrKuicvbadqo+Ur7nJW5g4F6q
BblvSC9rkgNB/5DyGMIvVoCNs9mPV9LegM9w1mwLa0ohLrGDBy2fxYUDIE5o4YfkgaCoasrl3cO9
P+mysyJCt3HPLVrjAE7hycE9XJtH/2gV0wRzm8Scocuf4ufzZzGQtCi03oYnz1K9fJHWh6bViIS0
8hw3ougQ9cHqQb0mflSBaDohDKqf+/KbI0+yTlcUO1GBIJXMypuOQwYRO7oGU9FpK8DhYyMnhUlm
KNWYv7T8RU9bf00uAMPWAc/heZ2AMMEi7ryWZeJNLl8yCLymNVnDUDo2GLt8oZZnNmfuSXK4FSTt
KwyM8X3Gn7xSbTFznt/i2+tiZ5dN3mbdJmFamW/y8HtyrsYs/UzrbSOn6fdTz0gl8X5imdXtIpYA
nrLayBG+6rmdgaP2B8piBun4UrxcUl6QmaN8GrWLkem4DRM/hxNskGSZiYosC4YrD6F279ExQHYS
0I+dSdWsmCJcwAAphwhf1odcipkTqzUx1m3fpF/LHVKUVRsf8rFSmLXdMMTUT8cz7fdbvjezXjE0
vCn7IFoyKd3EI2KeNBgSZj7FdzE7ADO4M7Sj7gC3JHfFmBX1AuH3feZbdEjZxRG7Zln1d2dd7Nwy
lcEg4pCxylOS4LFhS89rST63wmB/Y97r2FxJo5fJkPgkIPz4itJkSX+B8d97jkCLgPs/mHrFPu/K
mhT1tvHmCLIoMQurHNQRjs6z4Xb0GaMq/yweredgYtd3jBjBuuZM6OyNfD2lLAN7Qk74K0lQdqCW
gTgWls9RmcDxCyDp01aw0O4QLeZ/BpCUY3YB48dtcxsnmwHsMlrA8lKDczv4x1eKfl/RJu1xFJ0n
eKMRpT3H7VlLRXu3lnaydr3VksmJ6Kl2M0h39/IU3Ge81K3Dn2moz8E78TRujEtUqSaEOZluxipm
Kkp6tzgjk11eZBrbGutA4KW44b1SfEPaE+6UbwBcG+OOUxZbmKkBO/yLqXgPQI+an5qEZEcA8qR4
hKTnxPd5hOGdTqwUAssaTPMGhuxOTymjGPDRQWLlC1SG1b0qPn4WwSmrR3HYiGytjlXZ+5lctt8F
1bDOujolkW65Z0OB3+YqsKGxbUJ5Qp55Ppcj9X2o47uBpHqr50evsblZ4xl9aorLREENlLmgcBuc
zbQJ6+10k2cs6ZRpJYCW86lsNHUWayiDbcgu9KK9QPSbDsPiiR6tr0RZPm/NeVgy5MSr0jBSAD3B
ndHqiwA9tOuyJFCDW3VmKewYjB854+c3aIKH4sA9gMevE4e0ehUCzaH5Tdciz8zsNyI9sL6+jYT7
SCIWCQGTdNZkgJhTHpk62rXV026LShMpZcaJZCpavE/r9R2KZOh39uYJw7DjbjlDCuXlXEc491hy
cW6VvyAZVehIcvn71o/AortPUJH7b2VAdpbfTRrtLImHmu46k8yy4KKY8JUAQi5mE2YvoRMv67rL
gGM1Klz6dVaBoKS046RVVcCbji8JPtrPxqAeBTzitoYWtxFyFWN/QUudT45Y5LM5i7tY7B6fMo5M
VgyNZk70ptnvX99wKkRlJqXARb5Qao0FbMtA104IACxfGq5UCwpoIKP5/W8VkJXG3BIpabUVclbI
4eqf55Tfd/zMIdmTg/e2Jrnt06t/m3nXaxiXaAeqL2B+0EQu8oPgkXT1o9idLZYsG+NM4a/LndhM
sugD3R2xUlIjTj+yaD13edjuLSeR476kZf7f2csDbpNwmWjzls6WE+kXlgBZdRenFBsixb6pRzYE
L2NIAreeWF6wv7spWNI5Y4P8b9EWBt2z/SVaPVcdhJy5na81Z3KpgNsmhedAZ87qFYguHUCmyXMV
Yjdy+dDdU0zjIsZqzLQb2/+TVYXGaJyKS1LvADZbOu/83tGlLFjHQ0Jnqpw+tL9I/0yY9O/FGYOC
otNRCQyA7eBo+GY37paMqBeWMi+8SMN1DkJ8dnR3u412NAATXJ41zajs9Ek/1B5Of3rW4MT/4lew
FBcRg/Gs+XFcH53GkjyaF2Zk9SVpBxweTPG3Ty73NzfRhLzoJ5W60z3h4TlO0mmrB6IpokwXs0qc
8c45dLD6UNwxKJXbLe3aZky3/d7RkdXxkgRU43X0UIWkkZFu7yiVe6BOoJBXZyedsCZKm/oODcew
ZBfTW5/vOXW13pSHaAZ+nlkjRnlHHlSaIMF6fc8AfR/kob5bryQ3grSXuN+hKcFAD8boGkrT0JRu
sn0/dhsAphwuQ2bFLoUQD7WGW6Ra0npYsxCvfROJDgK+jcT081MKvgAniLUwBXg2zlJjLOSTglJY
hvPQnVU6hGqSOoFtZqwZCNqueg3fRyCIekdb0VmvGtLaDZciY0uc1H+lHy+QGqVQFjVsa5nCMUUe
VgnYsn41kVRdo2mtLL1ghruzmc2AHq9tAOI83ieTuIeJLD2I9m3GXynTh3Vn87aHStQXvSrsBa1j
hf6ZgtVvjSCY5vQPMgA6JPyisYksDy+xWkOi46r3ZogGGF7aSEGLTEd2gzY6y7gu0J5Tde7BtCnV
gyBkjEDG4T3QBg7SthDhcvFycebCDBExdgpLc4gV6OZD0jcHtgNQAHPDuSNqtaX4599fpHMecP8r
/5GRIJaBD5U7HEdBi46BHokvWn2V5mCF5hHgZ1SVIxZLb52+aRSXiTVqStslvoLYmO4I7Df+MFPq
AXqgH0Lfdzr8CMZXL9Zm/A5TYeSI2tg9TYDmgct77TLEFMy66dntRCVbOP1BqKRCP0jTuBcRFbWu
9JpGIU4PmTjgPuOim9+ppP0+F/jGV5vK06LNFvfMEcAr5X6oUEzUbkXKFMUKLA8+IwO0QtbSyuNI
yaNd1ma1aDmrQepLseXO/cI+tCT502hECIC5mhkpJQ7aq9TmMYflWN/4/kMhV8CqYBt9O6DO+9pS
Kx4pAwnKTSQfwEAOxL5BUIBHD8NR6w07Ku/1KcPamuYvzfD3hJfkyl7ZVTGv6jH7eSqHSfAobbxF
rzGyEmYOCRgU+HJe0lkcMvfxSj8yP9DzdvQnGsdGBNZFcwDvjbeQtmkLjP7W8k/xAUFyTatb36ba
jvHkQiyii2uKi6I8kZcnoBFufzJnUICxcePYULIlSWNrPcmwkDeRinYruy3+fcqFwXwMUdN+yrHW
U/AMXTOOrQG+fIIHYJxWMaWoD6QMiiLShEUxIsYj0VFoRzwPntGmI6wcD7Ff0KThG5PKi1L5cdtU
UUCWQv5AIzU2SaqkI71pEbHYIHw0pNZJngs4UXn00pnqbBGI4NqFd9A9kkRud51gvJCmyzENGhnR
ZJ49UEjXFEWJCzJTHMlM2ichJrkSaAOqKp+QRxu27eCU1n4AUxRmPwKPb2UtinMnZHfEzok4MQHF
wi4jBq+ims02zeLImlMK0Oz6mzplIWNSgRLkA00KdmrHnl8wjcZWKa5AiMs9PVJ4RJNb5XjWRLQv
9GqaXb0fAN0n074oe4UBq5XFIahlJb1btQFdeKG51uKKc/wGIDtC90ADhsbuBmZIISPv6ct5FudW
FAXXsuoceCWakaMoggJIGLEEl2zr9QJejZkqSPCYogMYuCDiUOQKyJR3iyo7n+GOPULJmn7uzHV0
P7rETPlrlEQG8DfTzCnzcfHSFUkiXQ3JyV9iwQqa1Da6XuBBFeXrUdT3YHEBJQoXpGHonHIMCmOX
G0YND7bWHjdDTw6E7mK7z6I2AxwdfjVBS8u6TG7p+nOyU6W30zAeoqTBNnWKsj83FBH5e9zy8kI0
RVRbvCCOqu9hIPMap7dzHYVg8uoT1FKCKeGMh/UJWURfjlbGsR3H6MQUp41vB2oQSUCltcUq3xHo
3/aeIejZ41BKcD1dBWuLSjET19znbeaNDt8EdFjyfSkGhlX1spGXtXLeVN8AwCKV3NN2oU2yWoLx
XjLzzvycXID7n2f1iahbxUTSrgUQMzwkD/BX1b+AxroyTG5R2CDbqmeE/t9QH4avpucIMQkTw1G0
yjTpHOTx10/2BacX4rHP3KBNZ8ZOqlQDg8qCe0S5KcAlDwtSb3fF04onTc5cpsxf+fV/tOK6YoIt
pJj7V9ubAVKHPud6fIIi+q+LtWlEYB+km2koPom2AeanZcXSQMwxaAtlhCZoA2KIXHBoV9J9TXGx
GUzmelo88wPNtnc0IbhYPao94t/yiIRXyhrySGomgQqvARVT0VqZyDoi40BwMK/w7PqrfjUsxEzo
GdP+sQhKWpCSf0wWSDl3TNNvU4OeD7fRpMwAKogZObZI7yXZEXQoNmBiF64zT9G8Eka4t68I2/xx
cE/RBSv4HoOqW/et00WshQmNZRRynGMaUkO+ohgczHgKrxof0/6m7jGKQFme+Wsyr9EfGmF/i/sS
XOTCSD6CWJBTCVOLHaJ5kpuql3ukHlGLlFefCbkOmOtg1x1M+64Wzzd3E+ilnolSr7XaCgbS5ycg
+iX9QbTnvOhKsvpWGpxbyXN8eGkeEzYtuLnaD4AoYKhqeLaXbY+Z5NTM5FNoB/iHupZZv0tXG6go
sXEs6yeSucB+xFw1gOmpfN/xxY9XD9iul+YeJatrFrWs7rI15J2E4rQGc3VmgnjB/rURB46hqakG
cjhH9DFLjcVIbFUZ/fAnMg/Ma5cIrW5Q+oqvsGcUkDCkagZ5o/7vw3KwHpqt5KlD3r4adSG0yUx6
GTytZMl6CIR7r0UoKZfIjBmJ2sILbvNUkZfKKIk73tbvACRxeW9KNRYmoz4xNKdMFl1YN3ydszvS
0h6JJpvbwFTPGy8iZoWiHUnkuXRtyvfon6wBuJUJeheWAVuqG4xi0tzgHBQnc1CwuBvwQLEioFdp
JpoVuNGSr0my3KQ5faTPeqGYxXxC1PQ1C5AupHVoK99Dx00y96tKs5gwbKCMTAWtPS/D1S0f0VK+
fOSALB/7p4P4Oq5dXnV+2jo5PUHFQ4EV1C9sDscfbOp3zjh+Sg8J72SzwDyuyR7CfaO+VOCHzBMR
U9IaTZAxapUMd0pGiJKsCzrGaY4tF1Kpb8iz/x8BRR0ZyiouF6Ik+KRZi3T+EyiSwRYTkJXu9hcr
4oGtOhNDjKQtDnc3hJ7sdt8UbkIh4UALabvACBqeAIcS16GtjlM5CGNyZoVr15BRx+gioB2wyIJs
cLDp9qcvjydbUK5/3iMF+cF9Tq2VXoCY96cX/1jiwQpxgKDy7EoaJ73d1tQ8+/pxjUrXWnB/zwq4
XwpyIg0pMV3Z+cW6zAcRHVbLesZnRlAsodUD++HLFj02Kral86Edid3JUepsQS0LcgUIJykEu0Ha
/6wlcvOv62YNlwEdWUeFW+hOvx/vC2Ef0ZgSB6apCd/Pa/YGYnI0eqD83eoAYxTGD9khhbL2M6em
ZUUU/mBIXWfPj2ZAoGxHKNFZcAZm0eljKG1JyYvm5ejVCaHWf/WYgU52otjo3CXmoeF8bsn0HfzB
kA2trHnvKMT34ZFzlGWh1QfD53cgqAIB46YYyR+kqj5NxNRJ6FIEG4yinvjxfHWONoea67xwKXA3
66ZzCCwDHLx/Y6GIoe2O8gWsQUr0WWQIsJhN+sZrsela16zJPKfQuQ9YPvnZk2/MX4jSsA6ermql
mWH8jkYLthiUSt2V0gjuJYk50yossU6PvLDzXVenhq8TSd9GEFzc8GkUOe1A6k2bfCy9Md94x/vN
gkO8JYqYMP+txH3sF8YqwwRHhSiLnEH7ELTZLILEHP+xusnyyX43Ib9tmrTk4z5aT0chFWgExHZh
9HWpNg9Ik7hztsCyeSZSMVjbf8KkF0mDPzp70D+MDKOBh0MJs/vLQu+70lliVVjBFa5PWenMfKGR
85FJyH5stZ6Dnw9ip36WvjPnZsgadR9FW+H9A5ZNNcSjiQHvZbuDUU0Ehzy/Nc+ErZLlz5l4NoS6
LgoVOcNsrrpksYQCjDI+fanV/o5wV39Z9iznnfadCe0z3t9tT8NZY8U9H9dQFM9ddTuAccJLFBRE
BhR0OeIDeozReQJ3EuPCAfK9HpRjptVuj80334w6+7H87yJJy9pGv2nIpKnvzvSYaUh6+OkPraO5
opydVGFUNzHOx0gLdfwbtObwa7p3L69rWoPrf+/QP93sHOOA5Sn/qrR77tEprk86lvy1FN5KoTsa
5+Y4PiW0u2RQizK4tUh+4PCDhBCBgju92B80VNiJJHJUh6UhNWm+6uNz9T2f4oas2pTVndck/kcZ
VKCxODCyjyP1js47dvDso5hA98hTGe06HTrEmP81fa6d1swIiMRMCi6TEvWq6y6blw+lU9b4CEUh
Lhem1GwvTBwpw3tOt4Xo5tExpD42yeX5FfK+WHxXkJw0aJhS7alqlcIP98MrejCvggD4scmdvdgV
R4j3QAyE1YyQneEGB0D5P0KL8aCUvisAOyDFbRPWF+am3nwaAIv24xd9rhz/V6RBCxs20yCZzcUi
UVGzWpyeJfrKAKYk1jqhbidzs7X6bv3OcbbkYr2asV8wFdPN2mUqwzNmVQhuOY5ldwJvtYaZ6Jkx
X/Nd1oOGN91NO7CMN+o3DXI8Px6JxMLKr17aGeOGYubKsRzfdQiSj1ES42tNBQNkgdkIC+FLK1Wb
fzSlwF79W2RtWMYTwMZc5revlMHmieZ8xBvPSB3a+Wj3okocc+GfKes/S1bDUVeBW/lpuDX9DGPw
we9LH2GxBsno+jeBmlXK+MUaXnxTymrSc1Sarpj8Dj0lA8YgO1uAtDVURL87JIYOmcUrGADH1uvM
SdWbNVvNZmsgIP4pVPW5AoioIOHLOmdJlsyJXnM95Co2YJWhBSyhJZYp+Zxtf5VuZz+/5ks8MdpH
uc1qaYFjOICU84pdryHG6VrDInLRh8mgRrjxVy62TsE9wFrK/tx3X3qhNPGZIk+ir6egLAYjaLKB
vHSOjnG7cs2hWRtqI/qSRwFJwsmInIAA/f9S7bpfn8hp+rWP3JbsLlpYp+0a7TA0j1iLMJU2lKvK
U3C5tksjxCDChNNMv8ScwUAqJMd1GLoMVIry+pzCFz05iD/nQS/WcM6v5xwr69aj57uvTuciIJFs
n7ztzOUDXwOWAQonywJneS81LgzbeIuLpK6rzXZuERLZo5LymYZqfoH/5eENA9KkEJnARvIZHkOJ
0rNzotnIs6nmVwCmLTi5KdryO+jIkLjziW1ryyef3WAjKJ3RnAIAVhPCAVfPfa/0BqznyCJL89Mn
u4dL8yoKerE7hWjppVA7n5Snov3WZzyB0wUQ6fZ4pOKYrENamCyPAQE/DapmcKUW3V1ugICQ1xmB
Egx2ZBzBE3xkmClCLAFJGwealW4qBmOzXkGPrGN+fjjlSgn85px9sJFGR9UlyEVA040w/Rlu2w7n
s8ioKu0u9d8xfcgD6uMBtZfy1mZpmHNBVdFFr0kJNKAnFGKpYwPqQb9BxjZmWMmWuq9TFJvsAkhN
qHPPQaeEZ7M04aFSN+jUoBvbGgwyf13Ng+g6VIW88PSH1acmICqldKfwMT6u/cF0TFMVe6qnAcBf
Pllmsa5vMp8LedSNZAzrMwj7URdtpiP7YFTljE7Mq0Mb2CfoP2x4LQDkQ39L+hXxLaRGJ1CE8Trd
IQTnr+eXIGX5sQr/7NXCqteHH+OOViKFXyfwQznzOB8Kl31yRPV3YGFlqWmGo7HDH7jUd0Lx31bk
zsmKFl533PzOZGieBQPaXNKX6Tef8ffrmBF7d5cz7VZd+AYrzaNyTUrFp7MqdzAg79GttxSObMx4
shwXVJha4w6xPhRMk1C6NC8IYqDO9dkFNsPtbBTSxSs3pqastoAc1116NF3qNFlDnsnTJIhuQu08
6m1Fp81fy0kp+gawE4G+CobhUTGELSpg0xEMz05UceOSi/gwh6QB/dKKi7/epWAVSuUHSfuSpn3/
nTzxwFapw1CCITI7QDIfte2o/KFzuCF4zVZ+u8yJQfVHNZ2DrsiA7S5QdonyhtwKMpQFOKi+OUKo
XlKlaWXkdY2y3+nCd/mOTTwjTdsM1VMtARq0rml+5gDMu1VSbeJv2RkYEtMKwyfNTPSWSKvVSXsZ
Rf+Qz03qEALnLFbZ3odv/TJKUJMfdgStPjdGtwW6MAJhMRdEHuCsRZKW4pXG5QB06R2giUbNcgkK
G/lOm4J1kvXEWagmHmLUoAhSh1UdQc+KfEGdOzrKHNVr4CPTdajsS7RCW6XCiUS/L4YzdNz2JsBB
i2lbctwi54l0/u6mS9c9dAheRt08+R2g0MzWqfxVmcVRig1yPE2rTTTu8TJsfXJsclHCT/UQ6O/Q
K7ux89XLnBQo1mncvGyqlVSpx7mj4kZ6BNM8Qumq/p+TsxAfd2n9qZja1tltc8PdLJtYSqWfliKW
en3iZLqoDSoGWhNW3NhcSZnAktK1Xk5slkQh5np1QaNe3Ljivwa00fRitr4eDT7GXYCe1ujhUIqe
5jAABWDz8m+SykzH1WgmTznJur4nrZeRUV77NBSy+ZMFJYDiJiQtnGj8jV9X9KCgNlIvLxfmXjrR
cHcN1nsSKSI2BScxf6Mt5VCIkEQoRJuR3f5Fmy1TjmVSHwc9rOy7phZHYDwMPmR0SgpxcbK4z1vJ
eOpJNbyYC0JovJJBjrl476ImKqvvwgIIcrTuhqqkJ0ocR9qXqy/TBkpJZuYrhHCXkjVFp5oo4oiw
IeapShepNFM3jMKwvJiN1ZqhMC5ivMH2BNmfWTvHW+oXN90zAwpaUP5THd25+akTMqWvQ5JB5cl4
5HKnMoj7NRVmiN7Ti9xOSpge2ZgfCnoGy6Y4jUmI2KfAPYTPTkfbQLReK371ACZqyQmPAQavSBk5
lzXmvXUGmyqgc4+tJTgmsO8Qi9LuyM8dpXBn+FDOvZnO1iFLTWMBItOoYWIB5ce2rL3M+b1qeD5P
cP4o3T5krgE4FFq9kORT7UduSKcuq4bSFR7pqgQgHrGktNR0T2zbC7ZPNVEgocEM6nugRQx8Rcby
sKvxXjH/9hdEOfZdS/VXd2e9AImYTQDALg3UsQIIWL808s564pvszo/BTMFG0lKsBjr0w8QsS8H5
Z+HRJFrK9mWRVmFmjJ6nYl6C1N2SjD5JSTMJjeELzKl8ljfOZNSGn/0sSZaDNH+nQend0tCZXo06
+35/7PftwQFGPP86Ld1O8i7HOUcEKFkBlxYZU8Zqw39Y2u0D7QE+pJJbVzS2NFUnU8u+dIfPM+Zh
xotZqU/wCIPg35V0DAAYOdUMkcWSEcfJmId8z9/KX0tb2phkoA4YDOQytvXbvcib9onxEET5hkoa
MezdpcKR8De7eXmYFrDUigzkCEM0TQ79xkirxnd7mAG6HixT51eYYg7NLdce7psfACB7kcJ2toiX
7A9S3LQ/CbrL3uaTO8w7HpnPHEVjz6OdOKqvcmqZ8BhOhl9aoRteXntv/EE8Ts2ml6cVEnYlOVR8
GLONXJzQnmeJWBQCgWMdqgwOUOe3SURXyHfVOzM2QZn41Yzb77wV5FONkktW9W1COpmS9hchELFX
G+laVkxMV+D97z2peYRm2EJW6ijLgrHGy7qa8WIxkbXe99hu/Hvp9Q1E5z12AiT9qGQD4z+Vio3d
FAoX9HzIEKkR/fxBr0z0LA1C4q8GJV2g0aHCIDzh1RNqtH20F/Lx+cIktipBB+Yu6Fe6kIqlVV0o
+qK1CAd11kIJRE+apycJoBx6/fb1xYyLv2owS/Haps3ODktQbHkJ2sfMHXQrzsjBS1RopIDyyezR
wNuGDkAXvvTAxQG+Hs5afbW2vdigvPg9ecLfyJGNoXH3lf6Y/2VrpMzJJ1O1ZOyXv0eeV0ese16L
4rY1CqymcIqABgQcr95UfiKdi+aYaVLvEFBx75bI6qbMI33cvkfASa+miqBLgC/oXO3+ZAfHxeqd
MU0HnojOPOr4itq0/3dn5Jya30Hmz5gwW1W+gAK5uhHyPfdIQUd7x+dumbXCQuERO7wnfTygQe1A
aHamEm97ZKpMvnTTtZ9TKcPSV040DoyS5YJcr8Nyj3HGOEv0fVEt5CekZL1WHQu6NVSNklkZ0dYQ
FIs+oyZ4Mj86CJYytWLL3kRRtereDgekOxj+3tSjgZjZguMBHys8CRIHhVDaCNQ5d30pD+2VDT3e
n4XzOGodPEHMliZoI3Z/SQ1ozilV76PDYReQ/uf4KPOd5OcB9LGyLHVTk/R62xkMAvuT1GqyOGFn
7NeXLZG3SrX6ll1znR4cXS/fesA4ehZaRSoO3RUIvQ/Qz0UD5wMBNWxmpupDg+/qQbbDvlCoS97p
SnCYfvWkkltOc7R1eT7+SdABDtBYmLcGwgZsK5daYIhD80k5lqvn8SsiNTDveWkPYPAxMQLi9+qg
L8arfj/qhw+fsR6nQvRSP1WWhr0Ecc76ht+L8FESFUcDooI4wi4iNCkOQ9JU+rLH0+FoxOZaFe/O
QvnEzvRrD1ZY5C4ckYy1uLj53y1TJd+U08nRDL37rpJ8xyU0t3H9K0/US8U6dNhY/dD3L+T7D1Fv
pcAMyxzZUOaPp5DiirdxwJUhTJMfALkGXHkUpAaGwJk/RCyG0pIn3GudtnprnrPlnXSh9VWnAjRB
3Y9h7WN/PbXq+RIw7sgv3Oe3a5IdF2SHo2pfnL3eBXSdHIT/nQ5uIbzzcIUZKRB/tHk43PrNU1LW
gWRttR1ewiXYcE3OkzBUPVpQpCYEWY5nOyq8GsgsFuy9F6raNcjueQ4NQYar4DCZHBw+W/+JmMYW
m+BQ3qR9M7ugIXZw1cj4F+9rcXTiUaqlwVNsWjQqfDwbGckhLhAaVq2+Sqz8UwIIL3TqQq0zDcEI
ew0CZVP4s1QCqF2hocr9fsSRQ0+7MS3RnUpdllJTRazVwblbarHkxmeEAlNzsiZziO90GLFsRv/I
PoQ3EYQiJ7Ekrvg36ddEfXcB7k7ZzLsF44FLrta99pDuHHgYCcavEsCRPVmqczREz3bw00Kk49/r
nV9t0sqETGF+ZMuMHB66nhE/RR87kQUI9Tdf4VB2f1NOY6mGQqBbebNTZMASFQ2Yue033rQHcpCP
SAuLsZCRTht2EjMbAyQthSzFG5Kxu9ETcOp5SBLQB0Uzn4hG43pCEl/Dt3T6xmd8YUqPkP4ZU4pz
Aw4RimH+OmqrtZbXP6FFyuQ4De/P7ct2XkXaMrn7UyYlDpwlqzBKisJn/ZJ67/9r8Y7zcRSuN85X
iXl21LavWTPSbZ8qgZIq1y/hOAqzuxnnictHxvFpH74ynKzmycVPa2V6gfBFv9J9lbyg9ZI3eecQ
Bouq4Y4z/wOK4TPfvRgLsxm25TKjRXVm+RVfryofXPm3Fl5PMtvDxgkgy2dEXUIgYYKEdvXa0JN0
ca7AR16lO+FKzfLxprUks+Rnt9Tu7eRELk8MLvP+uLDuJbLilYN5ahsqCSX5+LWFj5ektdTnJgFj
xBVsXxXvaEFTq5U+RDaJlzF2oAjAcwS4U65HelFnA0pHYAJ7quS838whgVYVTXmKfMxWafVOjqsN
u7I1/+WdozMMR6pZR+viSsX2iZsrEg954jRjCP9iIDk81h09nOJyPk1uXMbrNwsLW1imlLIM2dzw
DO2C418mk6aqmuqY0uR1r3VK6JrjZQQn0mmkZoUJPh8gzYyExmAUqZqrXfEyEjviYm7h5XUW/Fqq
xUhr4JOzd+kop+C2t+Ubkh1c8qzdrs4pSH9cxo2xXbGk5k9yL8Sq3JHsi8S63DxH2UFdhL4jozbl
uGatzfUWAiZoAj62qixEsZimKTOsZ2xpDG2WVbpkcpXIK5PzwSWZG2sIhz17qklcxdZxBZXt8M5S
tUBow/tzhkRRkwq/uRRJLDrcZPn1mjcxFxhizgWCh3Oo/WN+yl54hTSHquYq0SzbNCNj5Lqv8lHS
pX1pfAaKSzqBQ8WjPe7im5OG7F5FPMQjylbrrGXBCuWwMNtF8pVMHaYBuzSbmCkeP+ukC42i+ki7
G/NGXSMaLVQHrg8/jbj+kJtlZL65h94hYIRycIu3dL5/uQHbC+RF/GuJIfGbCuwzUw6j1YHjM9bb
rrxszX6dGniyAzE8XkaBrETCljIeP/4kMM0U+t26r4M/hplhbsNvpGBpO8RAfj42qT3/GVu2oEwV
aLyzctQrq43yq8XkKnshI3bEjv8MaPHEkRXuTk/fBAJXfedOAfDcyZ2GxtFXvylNcJclG0tlArPZ
Jsj4OrozknjTZQ8jMXpsH2EzF16FBZt8QIv9rFiVTybgkgSu3BgI+FYsthA6v86HCQkOhmFntP37
1QfmJgIp0trpa1bjzfRejP4PZmk2UF75YZarGHVob/Ek24K7bSz9wKc1Udjn3+IzZmeWm4t0Mw5Z
bU0DBpV6AShQkZEG0jKMKxE+Jod2Kc1yj+1SLw4Wp7RnI234mEvBLMBMOBqW8B9F8X+hEWLJbrma
+bEov2K6VtdBs+8BX5zWrFzMDB/NXuEVtI08d1CtHq+JIpEVjM9nacZ+uOD8psK8YK+tLQjuEx2Q
WCzkxY9YNSazrL383fTg0EzEb2IAY6AbFz2o6Z60lCaheaSQn3JNBX9Ef7asiu/rkh1HISwy4xYy
A5X/AMrObnNPvSHxmFA+oXCGqdEylcSC71lwoyszCCO6LGX5xevX/QmsG6VD97oHboGhQaMVZoIe
IQLIsJivtY83QxFW/R1xrhZ25Nx3r4SBNLuQ0KL4AkfFbnbROEzZ7BJL7XXTq0oCsMIIotPDrKjC
0k8FgypcBt2c/0w87RucNSq1xV8uXm2OwcOI7kak1xEBDaa5UZHLXtxJVBnZ/xW5PVKyaID+MANS
Vym4I810Moh28bQYmSFYOr2ViQPVg3zb11zAP9fYs5EhWSp29e/GFe7wUdMlTG3hxGK0pYVYiPr0
473TKlGJLAcjww005qnZP2TkJu/Ujo1iMVFbEq3FXwqRYUzMFua43L7rLSb1WuFUGpNxwfJ+52fi
4Fajz80w2cgpmGmHb6lpJiddl95doBPi4SZm83P4WcKqPv/arQhv2SWeketgHk0argSay10Ce1Pg
IpaxIJzGZOhJ5dRescb0VKHIubtgL3yyy/e4i62+MA7vQIiPFdVTSNsG5MNXyq6P+0mo8PBrp4Dw
8YGDolLGHvd1/qxfI0SVBrcN9ZYKfnHYeztYX3hM/I/17uesdFGoCiruP34Lkkdc3KXm55XFlkYJ
RZd4K9Yu8vf+yvbIhc6QfAKRr6JFHWU18sacdcmPFq1+lUxdc/RgJ03pPXj41Qer1fGbP5xKwsmH
i3JvxyMGAiEzxjcQKB59suV2T4s7Iqelb5MzIWaskPjQxX9CSHQGgcFfa9pedVwwHa2Mxp85jBaB
/SeF+13hLz1mlrYzmukSmY6p7+4i+mtcqXgyfOCgD0/Rzk1AVv6bm0Ta124jtg+K90uPv+22oaaj
QhbvP91So8FDo3e8mVVtga1S+C9BpsQbZyDCPPD11sMuInBUOmvxqQdPAK3HJKZhOOP/M4Jdknpn
wi9smfgm6Jb0AL6lrkPFUfSX4tSkUaGT9S5uOCXeHyijUt06h5fkeOKpEgkDxN1LILZ8+rTGhHMm
teyVnPMwNfZjKTC5aVlu+GMX2hxaRU9jC+YCmRCB8K6bfMLg9kHvo6fF+mCMsQEMe9yRhRdVodbc
o9WQhR4WgoMsXxXM8hF/0lIZLU3JvKmz/pI6tmHnselgmeGL7kDkEH+lGfF22dsOqKLGlKGe5+nW
T609APwRui+lP3RMHXOhBg1D2j3B5MdWh6FOrgex3Fg/YBy11UjqbMJCzgSO/lqEGlrHghJ/xDj+
E1zNprWsxXzukfIpTXT/gW/cNaUxhHZn8TdDO/mQoiJcLmY2PqSpUu66S67BLT0HJK/eKf5qDKCo
/1VqF/ROEYTavpbhRNX7g4PQ6tByj/9GtcN9uUeuzMMPOmdhRyo3v0ebFyisDfxUFYM58lNPrSbq
dt1D6/8u4RWt/ewebrkvf6JqAyY0kjKGQnIJl+4tE9m+mdJZTn+9w5wroO3RF//AAbrfm8OgfYbK
lBZRe0XV63DuN9CANEr2/7MHesG3BKfRgJrnf+UZcD5JyX8qZxZc6w01aq1hFZeWi2HTWKGRFao+
uMAzzHRpgNyAGBqCmHiFYMBerD/qulHyx3rSKeubncd/FUxW1gXRvGH6gyBauW5IXkKG7E7tgjU5
Mg6m7wzyXoypIrsAQn6uUK5Gm1rAZNCDYfxvArwx+mbFU/OUuJvhgm0YNCfo9jsCmOzdWb5e39ZE
WsrSd209646xCt8/5eBL6NMN0XHp4JV6pcu2Zmx5x/suOiHNB8bcyRsJ8Uxs+XsE9OG6xX8D7aB2
Iw7fEowD3g3ezyqtSjkPICNFvf5aYRvCdFgYTQSIq0a7Vmfz25ebobNXG3auCF00RVf28KLKYRzI
XtGD6GrVUjK5Gejkop+T/g1K+nxd+r0wamcO6CUvWVnTVgaTXpW9Ziy6VH1BniFCfmPjIIi9vBj+
kDbmw6Lel63B1tls0zLHZJnaOLQsRMFZarTkgx3jwXj15oPAtCG2pEtD7ma86oThuZ1zuCEr/f03
+egFCbYW6aEAF4TsCyLzPxQ++YxKsWihrk3aZCrTr/2jR6D9XH+O3N4+f2SrDl4HOovXw8VHLc1P
05yuH0ajRSOVECcRhAJYiOI6+pTUanBCcqeidxYPs/1YVx4v3jm37+ML//CraRRvv/0ZI1IuPOuc
pjG5nLrDd5jRxzswgf5BrhE9Za8PYR0eTL3p7LyS0tXCyWAd1wlzAcWKFlkB+A9oeOa719gd01gZ
kUdjkUIO484U7x0S2VvzPus48Cco3b+pKmJ45ufPrNGSULeg3bHA606asHlBgVOSbk2NHrwe+nVy
toxfOh0Ey1ZOFiiYgGdH5hqxcGXiaYk8bvfGHwqa4is86LlH8aeVNoGOCJRFfPWeQ8Q/X2GMYtO/
+kmwB4L9vtjvt+ZXUN3PwinVxZdwCb1Ft+vz3ajqIl5ZkkTs+//TMiSVM3c14udv7UV3S2S8g4gA
4IqHYU+55sSLQnRiH+lFHN8JQesBEht4KlTjpYu1wlR/1QAAWSOm9OTzrNaA5BPzG9ZIE4gXUXco
C3wdcPfKWIy2HvB5LlsNZs4CHKwet6LcVczvHVV7tQutlcgP1QNLLCKr0IFLy5l0CQU05N28Z2VF
49BfiDHZuGw/8+jhNmxTXXvNtzzwRxdqpHyNOjTeW9kZR0efSERo91E7ZZ00QMgcLwub7g6mnGEw
7gxohm9y+QYdmb7RHSOZi+LpCrmnyrExVeQ7xSCHCJLIB20zr/m6D4kJsZnQHciNiXbXLF5L4i/g
0+Gec2hmcY/hflSsXslDb0lQwhiCWjGpntCPH0iT67kU+ejTG7GtdLTK9YfcbvGfNwnqT0bsN88S
zfrzeheBnLldNIn9b/va8NBjXh0jgoOKRDHssjffCS3+Ifl8OVwy0hq0yGdwn4UJFvMb0n4h5tSw
MqH2n4i5SSZ/jZeQY02wKW0NP5Cw1BQoZ4PPSwyHlhCBsUhneIkA74Mxue0ziEmzp1R57j39V+08
E1W2VK7Dbv11ZQ11BX3Pk1g44AJAcPUTAMhVJPrP37HgknOUWo7oMY0Imz/rWWJAkQ+fmcupu8b1
0tQ36Tht59b8hdXJiX7ZGs97b1WMSw5NqetZLfsbLk0AJLEPJICMYI8AvwbGK1bJvZTP9D029WkH
mLbTKvNQRw9efAgCMzi+P6dKsPlgh8yekTFGRQTaBCH7pVY/JvOmqBpVbWLRZu2lW2Lcbm2+YE8Y
ayr2lMecHM8kBjXZP80aNrrbtABzOcDkRESN16DgLA4qQVqtUqM0oygdztIFlSBXbeoANlX4aZ/8
eIVEx4RK1i6rROZafpr1XFjyZCREsPcbP7qByC/5qrfgM7BNVweWmWCoFqPz3FbZhYt+wmRnIeF5
CjAjejkckKb6/AlZB8FVwDajNFaZdqF4gE7oUYGpj++sXbf8Lj8esRktMu28JjAGK+pruHNC2SSB
fYDmI5KVksU+6313POVtD7HCW+0u/t7shSbgxa9z4wv7YBH4mWX4bOheVVVt1ZpSYWSm3XC6Z9Az
oWzAbw4S5tu8ygqx/cOZPQ8EbjCqsJojpBwceVa0vlfabvc/lFMWA5YF5up/34RgO7QRPp4t3ZiC
br0mNka5+OTikU947Ve88Hp5YWL3U4MJSJ1qdICsrJveqBFpjRSxg6/wNfP30u5LZ/ZInwegI09j
g7IFsXpdhWDpCPVcukEVmDnpxFTR8oQ9t9GKVKLu7COL8oouBfcDUMVwmEPXA0NguUfdYxhV2n4A
V529nYaSbJTh4jSIGcebcLJNuklnTcNx8iAZZnBPDNVNAYt1G5veOIByZJn/0Ko6SdEVkFJJjEAG
IwFP+HgCZZC9vblUCJ7ZHmKAaFddW8iREil+Dz9boT6D7x7gywLKFot2lGBnftrdFKpmghwzVaIZ
RP0uQ8ib0FZbO1X+3Y2Rx/0REwdvaRRLXqTWp85Kz8dexnd95jW/OcWZuWa/gR0sttss5YhNp1Rf
aNL7W61Oy+mYGAjGwLGhA8hWfnLmkvhUhloi2KfM0nJeLiaf7VGgqY6+sQ6EA1CBVZ7Zmi1O9QpA
7Z/fncldrfl4CKNImOpHPWFUEVqLp8QTCpZU6+s85dpkpQzVwL/FYOl6hEgj4PG9hSqE07V7/JlZ
FEmoG1h9lewDKjQUGlKXUpud1n4p18AvG5dW6mdSt2ZKpBOxMj0rSQUfm3bNAeqgGxPYn4aEiFN5
i3wTox2M/8XLbbS5fDRr9lE1tsaw0rUdXRns+2vsgk8vccTKrklrx540BAsxZH4G6TgTAmYJnx1A
F74KVo1NJPlI00QpkqfmG7kM5+rI3NQ/ahpy8lJWtnAFtYaaWFzNFgEpVWYYLm+42hii5kykkR+D
91z1Wi0JZLS6lrktFt19IfYgjGXiZpmhMdJLSBgO7R3jzhrUO122bffDlftXXIJ0Z1Oe1H65xhDv
/mk8Rml/NNMOia6rJVwM56jHSd0s1GXrHrE2JDeLCJpXXSFY/zBMGgcQ4j55dJclgPdl1egagLrX
UfnQas8ykdU9XiYGKar/8CtzMoSHlBfNUe7ko1KuIMb1pAcKhCYuLdPa36FZ1V41RkEVQlhnDzdY
b4d0wjA9W9fmujuflciFS0aEJhg3oBbkzhaX4Zj9s0k0SW5ExceTKpqbVkL2pwFSogUswJ9q2uCS
wf3eqQ7fdfFaFxbqxJXHu1pyEp9/OMWSkS7Tc+RInrI9kjPvBy3pRCZJL5wRM5EcQL3ib8pfrtmZ
UqRxwCZULrR/C73cYjyD86yk3VgbWRI2yWS0VOkTiM8FYDOTZxNCGR8e9nfBJlesqsUt3bSppAjU
JoNN6jdhTGuLm/ecGVUaVScVinzQueg0wIeknewHQBLA5HjxUPcI+R/saD5PH56eTE+T19Yqq2i+
yxZZZHLPIA6lVuppz6D6am777tWDUG9pgeLxLgLeNzIqXJi5Aj4Q9NI775fmrMCkZIuSow06lHfb
Jj9i7cDznf7rd7bbbFSvoadGj11rhqRlNYpaxcCclciv8OridE1JWKv7gFy/u5BhfjrFemfMf5tQ
KL1MImhK94NUvYoBlFFKWW/k+boMr/y+K3OxGB501bPC4YSh8ovwK1FjNXGP0dUc6yd4zpKawiOL
vBMvdNdIbbp5tfUWiBKCUZVWOBxryv1TiOvzK/IkOxzIHBNkvm1tjn6SWxnhoC2+R10G4twf7AxV
FJK9lOFW597YKFMM2UI2G4cxkbpcMBkjUJb6XHTPDcaWWSEAFWnVxhDT/3JkO4tfdNtljZ3flRQB
7a7Xbn6TC5Ml6GODcnOQsRma8YkeGW56xQa5+b5WyYq9KCxD8TedQHC/7MUWroc/XuB2W3BWZhJE
t1dmNS3pUuYbTAcy/qtrN2fN+xKuuN27XSY3xrLXnHNip/x5JENO8SnEaYlHfVBrRNRLt2Q6+2jF
un2KFMapUApnRj4zI/9dCHb1WhyWNE2Jo5v5l88SJRjODnGLaLE4uoYc2z66gcDGnCOhTjf33gaw
U7R+heswl7u+N6WdO3biL7tIc1W1mN6ByFq45GqJp35NPtcucoWwf5PhYkLIE66bWEjXEt1pALvC
f2kNgjc6CDg1cwWp3RQvHXp7kCXK5falh6DSo4WXhINLIG8XqGyeKyg0jAmbmM8Gi2G1Dhu84Haj
dNVZCrEe0C8vCVqJN7BCcrQ0N81LopFrZkID2AYn09VMhm/JQzpnWjtmrCEuEme3S1BbbcceVV2X
nko+46cXSCm9Afgb0LOvn32ym1g4sOI2Urj7HYG7FD15ZofN471zW/tskkVmoBHdbfhpyhAXpoHu
Wuq/hBRwcCX/TBuXA7ReXQ6ybrs6NoDG0vB610Wn84eawBzd2I2JC5ScpYL8PvrslFv6HuggQhyS
lwdkR1gl+hY9HzPXu/niY+U7Fosg7JsGmTu3ECAC9iFm+7LBjTA3Slzh888N/SGvIbVvLkoRBdK6
L9sDn0G1qTAEf//xdzaoLVXMKuaFumRa0noJYnn/PELV/X2N0tBzPFQ8U5+AlfE1oC26PMue1Qy9
IIAWARLNZJDtaZeUB99dZ0sZo7zpzwkpU/xkxPP48Ic7PphKMRCYxh/9DuGv+CdGkQC6bK8M8Xb9
TsDSREaMZuMB7wRWUV6GhB9DGycmzr5LXdKNb736ti5ICUF1V6wMzK9OKh0RQpZdefc/ezCuvpTS
zXHLF8l7uroZljl/emq0flDdotbHFWh/NIguuGnwQhQ+t9zjCiP+6lqRE8EHuF17xefWZTs2UTth
1+ntTWutdyMnF+YuD/qY/mHg8uuaBKW9veGcrOcihjjykQ7+blFChQpMLcgQrOHZYBGfWFS9yJuP
0vbM01IZ+AyC6EEigr/Ckb9q0PhK0kJnnF/1H/14/VUiL36kgVV7wvSBsF1+XviPDmXYCjG9oALT
K9M8VSK+vQiDi3Ck/gKbAkjrKkj4Ct3RAryR5SGyn58ew45ScCHHbTfLDmEtwbn+FP+mzvmYAmT3
6IviqK24TIv6c8t6/lfZvU8SdX6WIFteJilKnpB5SxacFePZWNT67MATnINEZNvxfM/gnW8am0M2
irwXD/lAkO3xGjVptCUQTZtmWVpyQmsf4Us3q4r535eSygH61ePAs+ds03K3QJnNg5Ue9RQvK146
+RpDUkMRemsqHzsp9rsaBlpoWVSIyasJHUJU3cn95IASRwQ56QeamjLcac76ycOk8vSYCQmZnGzj
gXuFduR/tcuI1KsjdBQi6xTasXpRcmknsjxmFwasFY+a6ZGinoR5MtMuGpCvp5zXme5CfvrCSSvt
N9qgWzCmZfdZhZmbceBVCtaESg9Un5ZNbaaiPt5ZcV3p45RxLvT3ZKgbblI3TlI0glApdHI7rmLc
VWN80qoTeAlmJJOo8aJPHhc3glFw8y8OmLa5A5dehG91vWe7Dn5ytqDRRRgd6y0mjXgdJK/X1GS6
7TdrRi28G99HzLP313w6JOjwW8jFXtcfR42Vk2Z5Kg58MPrGXdYjQY/vZpZUfAlJdv8r4P2nQv3A
uFPyy3TFyJDugZghvb8d318aB+Jcxpc2d4Am96ymoMpSgnBKhqk8k6NhVnnfjv8FklAcK/Luht++
YsvhVGjZklHJfGCbhTcEVZSYbYMOo40qA4EP8qXEmE2lUjYFp4bAQp+oK85OBgMFBu6pmKzGwauD
riQELCdeiUhx1mUyU6TklsqQ/VJctC9VEuSwmDELOmEOw0MdnfpTJLg1wq43Yw0pns8fyVDtONXY
8iM5TUx4VaypnQFzgbzBwHW7IM3gOB9PdkUEB1cz3OlR6dxJn9t1oNwj5MfVSzG6kypWA4zaCGXh
aQzwwPBI5ULf3MRV7qkn+zeIjdP5f1yR7QE1eW04r+6G2TtogAOcCgxBXb3Coa5u1t+i7pLKoE48
72b+ErSSkDvf8jdHzjooXUr2MjB51ZRCVKUSNZj+qKD6zcv2U328JrKhg83V43R7PX2NsuzoW/qV
Xv7oK3X2gH0bh12ozjk1X2vILCGJXIBIzUYiB3VpvzmKNJRT1mtUdDAuc2NY1x3ZcUMqZlNPBK+w
vCZOkj0u7QQn+pq98w3NozVabXtvv43FYFxW040BFa11/KSMEb8Yg3rrA5KWtV0sHW3OWIVaYg9a
YaZB6sHLs/KfgE/zPrCnc2EqCdWUcqqq16ZnF4ZrNnrlyHTznN0au9WzXO8I/gGvD/nghTIZstsD
gb3hIQZaqETbbgY02TVmTrzamoD8j0aJww/HGwUxO5+s6g2OxjKCOgVarjyrizOIYq1UusjvKDCY
QJ6nqXivNOfwDdwzcWzGxCxBke9l2Gsc2yLp4nEZjkphCOHbnyfmHtR42Ykiq6tdhUVI451dLe5x
1COllZqk5EbOl7mB+7WrEC3y92zZFKmVYl5LXR8MkajM8b+UURmlsz1jjexBHY2RtkghF98jk697
ZJH2Ar+Xi4JPzk9NfK2zsy/c6fx7DTKboAfdCyRWTNaMSpDGsEC0sX3yO4jBebTDwwBqalkBaTI0
S57+5JLiWiILGcqTFApXjibQBLCtY/lG1+FjDy2ExMTqv+yN/ql0SJTn+nN4UzLQtqu1ujghKLbA
2DXwjqyxVZJPgCth3IYNY6iM4E3UpDP2ODxsC8qJO9cHCpV2iPFXPLgXjQ0iLPc5D660W5gFSOu3
4NgD166VXrGvq6pLSO9fOHBcqPaSOUwRganhVLzwysNhRRqFOiopOAMtDy8FZ9l9bvjSniwzv9Q6
1rJsC8W8KH/o4EP3mSdBsb5OWNC6vlHxW6tx8hpUkP45cMgFcLs/Qz0IhD4xIkK9FPb5YafgT5is
qKsJB4i+jE4VyauIgBk8xGu+K+hzegjp6b1N0jFSie2Cp2ELwR0YNGdyVdP8SNC1qTvmy0TMnXgS
3e0YfBdtTW3SMWOqrIuGJLaOv/hJf9NYSpy4rnu2IJNvzxlLBqsj3c+sjvoUJdIsfDEtknA8Fhgh
YtXpo9M7W9mJmyDVqL4FUXUGIf5bnL2K9XVBYQXOtbZaIjRfOeMWL4+ymQDjrsGJQK8Iem7U3h/m
n9S1mWffM8Jx6SSzUCeHMWVerQzFxR76N4R4TBNJEGRJmgN3dKtkIWf9BrkQWji7bNR1AVSw9JLG
ST/CfoVqfUQ825Nk50S9bkblOuCvC8a/OVwny5t48QJDRrPk5TzVILpJpApZRBtQQocdB+8+sgQ4
mMqacrP8YoA7zbFb+IWfXgpkKFaAvBbmilJNEXm6OPMeQN7nRnJXtBX4pF8lsbWYHTzNhrCIvSnT
xrOV5CgE03yTTMcRpWlEynewrNgM1i4QjjzXUOfx2QfB0vqFZxZlR5l+JIqhncwtv4sXqpj8Whir
+tNlFSobZ79fkJfMDNpmlXHL1ifYGdFDHGHYxFZPhyv/w1ooBwIAfHYSfi+vq9UGDek86su7fOSN
vNATKQfCW7DANMbmvzUfWATHi065ARhF+Tf4wyO1Z+PkMFPY6y6IJ4kDykK9+bFesiEdsDy4WC+G
gTIfUiiLyj2JgKeQCAedJtavJViH491pXmVxYmPvkeyX/x7YhTMcTzmFToLm7m7moagEFWI/5QaC
IzFbPQ0z9rV5vA02BOgoQFxMqPIFYknkCegxYqCP2+jfBQuwf/sjTm1ZqWZb0U6s3Jx01b2a3mNl
GV/GBqmAPVHgVLve+LS+5t/CEelOIf18pTtL0Y79gplRZI5iQJH+aqL47vCm7XWNcHzjsSkkT5JZ
cX6BozAGwiQn46cuIs6mfNEYtOFr/iyjOL9s2PEln6f1L72O1j0V7kBSt/aKAeH3y3bI2j21hmi1
eEWCIP5CWX+vGriA5H4gY0S22dc8ceP7hY/cHfFaP+pKKJ2zZEVeXQP5nUAvUpa9R6wPwZsYFlmo
QktLvA8NenBXYruZxY9SvikHUqhyVod0vCWxOMZ3uS+Bv+iYPb61cypy63z0MlN8e3zKqe1ygAMz
WjSb9PZAWbzCsIrVh+mS8Pewwwf6XADOqzki/Z6DMq74SJrU9yd2uDa2zI/s+UWGhTEqHdiZrgT2
IUNj0WYXyP9+QyB4uNt58C7MnGR89sc4avd0jPA+DUR8BHqo6w5H+AkNYbLAxANuQ5LnJdeKOJtI
LB5y8UEIAhUJPppI8Vr6KQ8U7VAXjPzqnWLNBYWimSyDQU6N3QUaYyg41Qpn82/G0LfaayLkKhnb
1VH9nMALkMT7Y7zadrtyXHX2DDYH8R+TnNXppOFqBvMX7Itl5LbCEhmyp5N/0AlKJ1ikE/M6yEbr
txf5YTyCw5m4He934iBwD+THEoTiZ5scsy6Z64F09UnhtCksA7SxkuyGSY2X1yUwSSXS90ASd1vz
QYv9n2C3bZVqOGro6S4i+8XFQbX/dsIxHiu7uKp2U27j2AvU+TZNrHcTiVeW6chqyMZHc0eTKCeU
6DzMnQbTrTKIQg663CgEC9iLxZnpqap2bI/VkvEkF5cQHDpgUeyA54B3ExT9XdBwFciN4KH3lmPc
VMGDTyuCiTv9IlPwzZQXba4Tq5pF+YHxuP5G6ijbLoEpcyaLh1rQxZ635AoyL7tTePNOpf/phalf
dbhj3j/B3qPVPpnocLoc9hfVesI0o21AUKH2dwJ6n4wXIgIzX+z7/vSuwhx0YAuE4Xg2/udjTASa
/NAoK5N81V+OisD/6bI0PCT+gvEq/iYlg+oDby7RcwzDHRHP3+FBD4qFTuXs+1lyvHNU/m7/zuC5
xgiHrWm2nuNDMObASvco6zY0S8fOqVUsyP2IIs4bNbnOMP5ABTaZ/N3YkTt99SflxE298lFLR7LO
us+nRuHIppVFTtnCawDLOXn6oGmS3eGvcndrATB4//7lXGUk2q2/tV8HWgPyGKfEXIKiDMB2M2Xv
90iO0YNAUwT6a7ELE1R7tbKn2D8eMrv6EcmFjCfEw1tigIYVEIMYv6l5URdyCQsxdNgIUlwQjwEo
8cOzF9sq2RILup0GXQMR9/HsutJXeQmgYGdSObfNa63ETrWevr+ag3OYMlicQsj4rUAFByz+1G8P
D4p8SCzP7SYrWt+za5zb+H9sLYUUCarXYYtAQMbNsROaupX6nrK80R66PECPWYckGKNKSMSzwF02
AQRHAhc+9Ww52eKMaT3/Qbjv4/bZymhZIOGJhxvv+vurjgryxJQ711aOJ8XyxJl0RmvZssawik5H
PN4YR+LKE0PueYb4b1xN5nSHA6RfgjS8dNBbJrpw+jBGpA9KEiZOMUUYa6MoRjCFVYC9dlRxCCP8
U96NZtp0DKHRnuFkLioDkh4On+bAczc8TOj3FGYbEhe0O6/xtHXoskxz2jvMnihJSUPsOW0Gk7ST
qcsKWH6eU/Ru9xSQcAOVkAz4qKZHqCKvjqAeBbNcemx/lMUNzIAo06s53RizpQEVE4ygKSlQrIRZ
0oy9A19574T5ZgfCd2nwuLOPCMMbRPP88Dq0Zj/kv2ekeqbWlBkQhqhCAg0stSrMkF5pxGBiaB2t
w57F9CKTYWvnP6ES5UMTXfKDgycTJrw/6RBeQ5XtrZ6SXr3mZLu/5oRnYiYE84tpbRUMr8V6Y/Kf
pPLoaT1s4ttgqoXs1rytKim/b6+AIX/qdlRQnvJz4Q62an4wweinLiGoSg9BIyioilkFJ0QK2GsX
/jEZ4bEnEBro1PGF414L9g2fgTz9h9SIsda5IspTnuuc+V4txFfHSshvdA7H/uhepm1hP6NN+VRH
Md4UulqLjqIKEHqH3m8mb4mwDU8xheP3qNloARsIf5/aDaVFb8cEMjJncPvnZ6vPrK6KluRkLDnW
dTbNtS6bF/NbGaXCQH+iyo+fkZwYFvQ01rf05KhFM3TbrX+HtSlEBgblRbx1YxRZBLjumxUibROr
mBkB82gqrSWTEqIx8Zcwt0Ail47UD0zIj9OE4gjMkkQM7WDdh7OVshy5FG6YIprFDfTmNmmFRyxp
gATPXBBv0QYuTWWqzFecAxz40hO985RsP7Tlr7dw384M7iEzBMBQOGd+gZMuh9HHo7aDFdAnoyF+
sIvi0nTNqPTwsYejhIs7mplUAv0n6fN56rdO7xprCiF58cxyIT+3+qv/xz5fH7AQvIIWX+u7jX/k
uowD3LzaXgUPUlJgPjQIoBAN1cwoSqAGJSTFAjUYVyshQMGgMeQRplFang6gHMyFefKLiqrwsOw5
qgtgSTYDUw8W3xy6Uah6YOMsuWofD1LMmsUow7twJ6WzTGbXV3dpxXa6vaw1BodD3c25DWmJ2kJb
nS4HU8fsq1RngBeVyADyte0grQsmlORTVFEk06gO2K3x1k1CHX1ImI8/2v+k2oPOyChDVS6k9Tw8
GEq3AXjfyMH0QfyYiSd9X26z/JPAr03W5NPcTL8Z/knU35ZYbxKYS07TTfqE2nbV557+EVplt2Ds
5VXyfdk4szbXKGH31jVk1dnYhHWqJBBvRmTXlGYkd0VT5rhG87dXlWhWLgFibE7nT/CnyB/NBHUA
47nazOROyGtLlMqzOpDHwyL4ORPqgFSPlaJFn9a8JQU6TlSOjdF4h34EajVnpjbvETWv536yvubS
2D/yUV4KPhNRh9cm50uWtYWRcqCEH4HalpmPsOUh5tLDc2zAeNXnhWrRMzqet6lWlxz/2+JTlYEa
S9/Xg+2g/TOgInWgI6Mzyu68rN7DNkwHOOjAI4IKfXZG7a+zAO0d0ajuxN1Om71/U+Ghpdw3Kz+k
jXGblaB0EByocZ/sxBjvgDQ+AajdniFMhgzz9KYCqUD84vRtJ7HEBHYjfu2Qk/0/qs/m1+V8eRC/
kOD6HSlzZ6YxZ6Z/OhGpW4imSCxZioLAbUjHWjKa7E/JnuL7fKAzbyz3aNGf/sAizz6Tcf/RP+52
Zpg4p2HFY5dF76xWMI6oAPIrFB0kSIKsnN3uZp+LclauETbZ6A9bvn+FVsXSQmRiRcKsADwZ5OwL
JDo5YrtMXek8ty8hPKJgujpSP78v9DdimhSuHQJ7uVeVPY8kp7pxJaPZx8xCCoes6Alfo5+vYcJx
aMnyTrfmTX2nMsHSkTuV8+wneeEd4EXChQCFDVzq4pyhtzr6Vw82AlcEaeZfwPYC6rTyroacnU7E
yYjA1C9n9w6YGh4MQ3bDTPUmCUywCV26uhcwNTuAMt+vnJjXaNFT6V6IwkXpflsRTY6KFq8EwjdQ
IRoWvvPyQ9aVlfdFJ+6lFMVGultSKv+YYQ5QSn/8/wUC8LAj++DaXydNTJtBIwgLBJrpVT3L4Ajj
SNwd/YkqVCDcgEv54ygfkqe4wONlElxxBUTmNuFHKMvH8e8Jdzj0kMgbX30CLTzZoLd22SldQPrO
LlAUkBhDDjJeFUcX966f2VJB1OjkpTJ2Z7mtbQUMP1syA2rpoLjxsjy5rdw7H71J3n1f5rEE9bab
okPt5wXfxq55milU5hpcJmnqqsAWjFS6NxdDhxgXQb44+S0TNQld4kBAk4NrCb+TZ6uDT8ClUTK7
qTTc4oZ5guDs28pLRCpZYPRCU/+9dNgx7+Zj48UGYUKAnrhStBSpXRqSCAZU+5LQxLqbCYq8hdqQ
mqCZIrF+hlYBpIuuCcsmRySfy1m5Zwkwt2yh1hlNN4/DKoQgjiRWZqheuz4HLL6A3bSL41DlNDpn
ytYwxxK8TGky/NLj/zubxL7cBcasumiPiOEGTo2Q9H25gTsRzzWUgeY8Q88xcHPXQzVP/eCvjh/q
2Kc8UR0svSt6lzoUU4ZrMZCbf6AT6TfuyBxS6T/ToetaiiD1kB8Uu/dfFoJjdgf/Bh2Bcvq9ncqc
3Sxgzbz2uTYhu1VBQo4DkGzsZBcpf5pSgU5x7Fob2DEJmGXb1d11Qar6SV9PnMJwxvEks30loVGe
/zvXxIRIq4nb9pxfu0jL7AFgg4wrwajFEcLpN/ch/u0iCnEWz7PXlRbU6zTDtIuu+tBgPhsD53Qz
KJrA2o1XpP3XgTeXnY4vr01uWB6wvsG1D52vWguevv+gxns48hya7RFBKssuv19kjV52E9XhMLcB
Zk49nPGaUIpzllFD264ekzsU4lhlMj2p7lUhtN5cUDfJm3jsupUNqYeeBRC5CmD+JQ4rPU/MoKqe
1DHl3VFCDBjTIz9/6Mtk7VlegvN1oDCkmMukjCNtYQWGV20tlz87/tmqHroBgWD2HttI895Lldm/
NlKB1kA4FjbLv/Hi/eD3U4gtjlgz2SKPkKynpaOB0e19s1xgnE068LwoN64y6NLzcQyiBA3hvRCN
ZzSc9YHIQURE0Mxc7WTVX8ZBvnFFbJ5pLwJoVsp+F+t8AJSF/GnDTrmk9o1/kIs9NCSyfMA/ZdQr
XeyLZa6ZdeVb037m0uhYp4YEP5EJarLuyE0btYmRO+0qApv8lzCsZFk0zp7msdOgiDAPHdPHFG7t
3Bgf5g695fcAzXsGgvn1CMjgVSjc6qONBjT8NZyCXuFR6TG6yBLMdwyBSgs2+57oV6ZnitT/wg0V
6K/u3CKyrXUaZT3bQ1/Wj18XnaGIlQE34rESQ6g4Iw4yCXmrLor4cKAm5jiox38DzBHBDLhoRRKt
HbDiQcLHDd+r3RhwTR3aoAimjK/V1o8F/QxV8dgk4bqSayRfhmlzMweddIgXEL/RfkFViFajFd8n
XA268Yq8149T3oPtQFXUknCHZj0yWR380h36iCcR73xn2nnNjkAy3/pId96a9BJ0wdCMuacWewTq
skkrfTEJb50iDogy515diCXmet5gY7cZF1sZoyzZxMAAedmM324LJd9apFu7AUvB+k1/9ZKXAFTv
GDULWIECNNzsE+XTm/Mz9Q/DhzWl3xt1R6pzC+iG/v/TT3Eby1N1/83nLyswJ05l804NGLfK1nSr
UvKZ1zQM9jxBlPzJwPewo7GPi3ck4GoJpw6wFXX6TwHTBbnAuB+07p9EwDpgBL2IqGcpMZMhkkS6
OSwniiPaf9C2I/9avF0+MHlOwzQ8le2M4rUGoTJHLxWpc/KTWlQjblKw7B5vipu9wQMlzRODO0CU
Wfh6PHJ+vcpt4Pnx0vck2n1Zq5t2MKbfqznUpkm94zT3t1MrEMSrYouZ2BTAkgTk6ZLuM8AzMiMc
/1AS6VY++50rBMuxUzyzDMnX2p0DHuWIop7iEb8aQUhZ5axNqJdM3AsbNzXy/u8sbk4SBGb6oBL0
93NrZEzJkOr4vBDAFxjQQCR9VQH8HYDCnzqcmDlJ4Fvwio66HcDIn9rHIZ/vlrtK1CS5x0mxzKt3
JWDCeIZdZsbJhEZCS8v8uqXJJHsep8DB0HvJbnuc2uZG+Vv3i40Lw9COmbvDXjKB7oelG2yJLhZO
AUHx4veIMZo4jN2+hDfyrD60mUVqIGByrthKxRfWCMYP04bD9yy0DBoBS7jA3A4JzDAKT0s4RnJ1
KGHJ8MONATPCaFzblIXkV5rZbQxHpKGMdYgPmkKwrB4zrXusffgvwR14uuNH+1JJ1HH5LTJQQwpf
zUiYAbD+OAPFEeLuKlb7hXl4zXrMErVKkt2k2fVmwjBQv3nR6aH8PtctjnE9uXWmLNmQ2VYYep5L
/+l4iGAP6PjD5O3MISfx/PWo88xk90new5zh1cpC190ii0/Sjx2XkqOTNqaT0F/bvAjMflen4sqz
iMMtFwdqRKSS4puwsxyahPWXXB1jond/uVu39YuQID0DQAP+zM1z72OL6RkX8jR1zBMe5v0jmQP7
Rd7XMxfdaVkzRmheDy6l3Ak1+T7BCn8E0IJcQnsNuf8JiZTW6GW1Cog2JgSR/3h7HgX0gRz0D++Y
Uj9QzCbd8VFBjGbN0/YfssOzwaRaRPuRIl0G5WboK96ntro6RX6zjg0l/3IKe/9SM6RaMFu5RP8Q
9umpuKgosdeu6vGqJL5oiNeJPvx5EGTkzGoKpS1+0RAnzF2wtUM2Ue8pOlvVLS83aXa7QltqatPy
NxtsDOll0VF4Ti7SIW4OC9svLPxlDmdvoGlRH1wrVM+1lbgbkXQJQBtIFFYzi/1s71ThACzwHqQ1
j9TNO2Jn/MYIfPmlNmPAPtswgMsdYGPIejv5ywrNAtaEleGE//Vl68ZCZG8Xlm1X/l9was1O451v
LF5goCnso22iztMpIx4JAJtqQ4uEgKeZnyFk1hfLFRPaXkwAGVR5KDrkHnKfUIbzjNKeDlqhTLUL
p5FEe0SvON1R2xVoZ+r30C1soquPAqCJcXeuIGCPVXDz1dwsXnUdl9A7EsnHfJWTt/UJAygOzctE
eZX7uv2EJLBySr/FQfRNB0zHGAIc6EFqRB2YkGwbBHZIAERtgH4yAl3oRXq57nopuCgszvPASsjo
OT72SEl9loQAMdNnJvb71dV0bq2rTWdUcud3jdWVjZnoajgftuwVlcuzUU53Z8NypryK4pq62QZY
b1J9hMIPyIQIDjoriR9UWJOeo+BNo1bvt4ntD1451vDJOcKSgnS4ataut3guPwmfcgNkmPw6FoXz
sxE6Zi/mEhiN20mXktRO/ANVC3+quocev2NgvwDsm0UYkUkDizFOscBZS3tTdoj0/1V8cc6zyb0o
ewf6hlh7PXkTMMUrIWw8TAWftzbEXTsZLAZYE6GjEAfEAIztd9YklFTD0BZbhRnJYijQE1HBTfYZ
2dl+F+py/15Zl31aBJfJabuSIvK3uk2eGXYDs64K1uQBIP1MUBXbevl4qXjDDPcgsNc6yX/wkN9V
T3rbmCGKe0uIhdUCp+kUpoHz9fpZEX4T4hSoX0KdY/kYl63iaWUpsASuZtQnPXmWAyttfR7r7y85
qdjbRDe+oXvzYjQN8gEvYVoiAE0zLviDAbMACLHKyek7XRaxGXeWYb6wqnvnIuaYe3BsvcNPoaqe
XDv8zroSQTqoC3gFYYRReWluEUVVqdBQp9+SoKwBX0virJDpYZMiTYc74TSteGDCzYf2ei1UqK4h
hS8U+9RgJjStt+ndKkC2RwuMRQwqYOusu1eh5CZhcglB4/TzvdwM4laafOuy/CrRSa5eHnnGiP9O
Y989h/GQ3+ZtlgvQLEm+CFn49xoZAWJ9DUj05dLVJT29iVjeBbq+eW58+UR6Sr638sO8f3DBe2Zs
7T4EiW4JRNd2KiMJ9FOY6y7ahGU0bXp0gXMakw0/149U/b8OxcuuriY1fSDlWB09zAtLcWuDFj4v
ZxlxQJrSerCtzOyvvVcyV0h5jkuMBl2e6fLGY6F9GZ6l8nqAjBSv9ogqxmhVoCvfnzCO3AugR90s
KTBALecpduVv9wT8qavW33JUyBTQN/HVfYilkNptaLG7b+c+7l6dDrJswtdM7qjXpHxaHjFpQfCG
2M72KfKaNd1aT1qeZCAen3ZhbNNTAhO71l6Mv3VA0EWb58moZ4vLMxgaiMobdAZ4RJAgfQ5GHRZU
+Qod+8LdzLuEMfO0OXCz6fWxDSFEP6HzfhFUS8dRe9jNxWC8QVOcO4FSjOGoI3gS4bGFnFx5XwHM
/ha4ka8AdTWcsDhH/PWEM/GpYNaXDmVFc81Al7M1asxKnu3JxuoBR/q63y4x68/GpnG+KKgtj1NU
WF1/ZGMLL4u9yF3KOZnLkNdUXC42Yf7KuwFLaf3x/IZv2M5jrvMjDlFOpC22ikc+sIvDSh4aM9/C
0hTM57cOhvR2JAD3ANE9duHPogQIGa2bw0EI9h+LoK3Prlzf1tyaNsHIDNgR9TfY1sz2wEPdtjfS
e9E3DdPka4ITfqeI1C4q/wEXr4wZzc9EsCthc9Cetdj3x/L+RbdBkCPxEgkQWpUW4nzPlkIw4PtM
THoz1aj9AimRfSattgjODQBOJqQUcly/SXDjX7jmxXLN5Vh89OqkJ7zHNc8v5zjvt7GxMsmiDlzq
hWDTt+EQiCUQlggtUSqPSd6/Yp+V8jp2w0gkpiIsjeWvOxspT3UFQL6fOm/pAcon/Dq1EiTnzsiS
RaLWYLgdGfE9sj72siuJRCqDZiEFZ2HtB34L+a3hQb36f6U+zjuefMBYWMATClwfzLZtZWKMsCmN
SzVI+xacKh9TEfr0vGI9RLy7eKpDFJF/aMKkqU/B2Y9KyOlkGw6SnGD3Ku6Xq11wBactxO6FnoWn
anNuFeQgQOrDhRqHck2Le25E0bGV67VccMCGc7rL2oQpq8HmBBNJcfW3dEBBnq5lEcESTAm1oV3b
Ay/FGbFpWQ2oxGFgNg6DzzjYoT5s9n4uxMFWWKwUpo/Ct375SBAaUL503ztGPaaYHsLGOb3NM+AB
EcUjE5B92pNbH/7wFDBPZdUtW2Lob/qO/F0vEuznHPAHD3JBIiiWOyGoFJDexI8TSsBT4/myD1l5
fPw1f8qiDJ6fTK441KNz0p9wIByScevH2rRIWxDzk171DE96+ei4/YTxG+lVhoMI0PVzfDtyaK99
/bLY6F3aFRrTu+q2h3IIFJCEVEH1KDnNbU7uoQ3VHDbusWdEWJXXkw90E22k5yqfm/HzwnIYd9dw
l6uF4WXNvbGW398KGCO8sk7EoL4BhQidl0F8CBuNgmWttI5xVGyfHSj/w4xKTb7GUK4Fp62XU4an
sGUOefcGmfN6iDk9aJHIB5JSSuSE3PPXEKkOiX2yfS6/Zblf2l8SQUAQRQm7jegYg1LHZJZGyNUM
xuWygkSptU8tI0XUh6YQgoncceUitCthdcrOEOUgcZ0B5BtSqp8jayxDTXD+t1LskO6i4FJuDJ3z
aR2zjXTIQ31Bk33pooFwAj2Y6AGhOJHUeAgtohExrZWTYlPXP7A6Vh8d/8IiOYbgzTrfj3qJ/z3B
x+MjvpGqYAlF+pPkNIJlG6Y6ZTYV25OVYj9g/XONHBwEweWPjcFfRFW/yxjuHPb2e9o6CPJu3Hh2
OWHTDzzGF+jGEs1sy1nTixE5i3ZcWPFNiOzloUW63Q3AageiUUclyUF2ydAQcDZMu/uFhscv0d6e
0NbMpHO4eUI8oOLKSsEXCvWLlJCWGIY4Lq6HiJ4UYJo2J+6zueqvq3yhoE/R6NWsgnb/HXpFC6E1
pw40mF1nOVM1++vZbXehVV7Mj0OnC268biyN0e7oyu0BRwKs4Mv6kUPMFaae3iz+QtxfsJOK56dG
A2ylXH0/OjCDHd8UxrDUUhoJWxsPEQx/zSejl7xH4GlEnASUngtilsTwhYlbygi7nk/ot46/oG+p
NW4Ty9vUjecdEtk8NC57eTWYzWI8g6MXpgIK4p/KZlLoi0dFCXsKj/fzEOobMs8hPLEaz6gk/Yhq
ysap5NzAnDsFGnAB5yjvr/4mt8rf8fYWoMc4fJOonQCMKIktRkq1YoqdB2oCThRYnwsTVlEglCcE
0vm3dkrvB8rvu5OYx2eawB9p+Ekh1Gxp3VbwSzvOlE9vKBA20oHLG1FqO1RFp7Bh0xUADg18Ne+D
Hdxcb0p3hP6gKhU1q2nh5lhAa1NYn5YAX4knq8OhUzvFTBCHfDIpjTXc+TpTRXK1hO4PX0054HOB
U+PCOyHJzY4KRBWXVmsBAMRsWz51v2wh1XhTWz52LVAD9NQyX0vClNj1ByA966cEaLOHZC+z6tPp
Wu02qmxoo2OmZkeCo0RW33NmCVtA2RuwZQltgCm7Dyg24/EdwR/TNg03PR1add0Q37Uk4JXoJb2g
Hkcoy6ua8ZzbsDoEetjxZarHeDBQWJwR9EMU7VAthiCIloh3ncuNdtYFpoKAzXFEqIOizAeAhmJo
Jk4qd/+Ihw0xp51QOnkZX19g0z9jaPM7FRSEFojklvtX6NXAZ4V2F12uUskkzPWvYS8qACVovGUT
aaFtAUQj3XbGAjwCUcg+YVQf6mWP2nsljvE798VSnp6l1v9PH+QQ3lfWsfBYeCgffcMhYy/TRGvw
92yCLbloqRgFX/oYN5o49AMPc5dMwC+ndVBKQ6sSaRBmgrO41dpYUdh6+AJmZIiPuHnjRWrtuIR3
GEn2BDOyAIC4s+/lbY/A93kdKOI76HzeadluxE8GnviVSu2cdv/VmtbQ1V1yZ9jv7nfTY67E/cxL
K46FgHaS84APN54KfByip3deAk5vD+Q47q2ZAq68TV018YWxu9nNTzkLFJ1vu6XlDZjwG1JxC8kB
rMdIlMfJUevRpb8oCm0Fwe1Ofg3kH9U9ibqumXmTQzj/FOoEbIehsVAEOtMMCGHQmwDKzYqJqbVQ
OjC/4Sr83lfhie7a/SRphp3OdfS7CGeizEMbE8jCrCBz0ri7Zk6hQxULC8OzUOwPDI2LDhd2eSk5
rNK2Wj7A3VSVqyng4A8B+37nZzO29BwNRa1Xbppw1qEgDbt3SJ2UnZfH0ZyW6QJS0RmYbeWpsiDy
ackpyzAdtiAaaM09Yu4YrQ6G9uxUh2GLduR62lUGiWt6ptIMad1dOFVjkHgZWTiNs0AYA+dqObNZ
z+15qFAThRY8W5ZzaDdNH37oZ+U8GM7FDT9pjtA8KU8pWmdCkXBg5cqNinuAMjocrXUHXbrLx45W
Y6cmTZ5ZgEdF3tZF9lwcmxZhfqwKYLVRbuXHn40gMiAmvmKoCQ8rnFTOYSDEva5tdYZZCnCZcXo2
4Gx0gW2jf+wDqYSus17uWRDCM1E5RGFyVWnzUNjJJpKEQSAloOBxTxAmASPb8iCe7cnaXHIEIBSY
mZYC0vbDoUerhyeXWvLnAycSZWJeDZen7Yu3H7NuiWKAGCFO18hek8lcgWv7eE5R0UR+8FrrnD87
NgFVrw3638xdJ5WkPLPX3XWHrsELX4juP9ejZLnlpWs1ONNUR2cEgqS7ki6y2n1nVgfY/fcjqECa
yn0/bEhXDgSBiA9+ThxJTtYyUPAKMtVV8QEkC/TzkA36TVNvZHn9kcgwq25GWZ4PGJFYEbqX8brY
SyHyX9Wpl68vvnmQBwaIKTkD8F2azV8jFntDPaySNypDRe3Q+FSNIHFIqq39cNK46QHBZksMCC47
6H+uOmy90ClUSi8fNFD30SECal19M4CwaQkrMOyB8btp7JpMuQc1DtgWYoaRgvi15suOAauURo0F
OQr3BjLvG7A6UW2UcUGkjtfKJ3mU59t1UrcFUI5Wj4gXNyYI2TzcQ0vMfRWQjozT6h2MeRyik3O/
Lz1LAFskbZNUuhoJ7JP23MwrRP25TuulR+cdzACA/1u+/94CSiADwRAugwygWE1JBO/JK/TqdEnL
l7xyhu3DJ8u5LBi+USTShGNYgOm0Xg0RjHOeLwjFrBoTOGKummdmxps2j2EfGiToACT8To5h4ELz
iuQ/nL3nO7i5HB57/BwPw1k0szwB/XNWYPVHv6jDmEpQ6LvOkuEdBqQI5fGW6nKiuJiF+WSYEzNg
yC8UrBisPJo5+Kn1rCzhQsvHwGGi/kXmUgCu9gcLzjazEmrJqacwd8Nfnp8r9ZlaaRTYLFlomxpe
c8aOZFSlIoWVk7UGNVgllDzKgayt4OLb21EAs4gp2pLyGxZ9EJGVmoAbbhtK8QNJsKqjOP34wQCg
NG5t6nwZRGgQDnM/FWDW6rMwJibm+vxOrqDWB3rlLE2m0ecONeEzFNYRAUlo55rIjyW1rpubXpX4
Jyy8APTQ9ZngmfsSREIyN4NaGMo+2I4jAAxHHRBQW2bimZrHwbwgH+xfcibyGQiE6/CZLwRE/fHO
EsxCli3JAGQFafg8VRBggavuhut+5Fitkd75wyNpAtgvEcywzGx1rdQ/2cPauiGZodBMXPBmAxQY
aBZncZCCNd/oNTRZ/FY+8ireROrGURRz2AquFFxwWLBFfOO/AJCo4UsRjtZr8Ib4fJcUEH9RfByC
39+wQwXyE+E/J6yjgsSmqvdDKKciZLURotJ2ZdbUidzY+vKbCndaACFTWZXBXIeZKmw33KA0GoIF
IivFhtsfQBcktouRzvOFO9Na0ZG9dMkR+xKMalwvHvWu8a7JDg5hh8ib7nc3wjWVpQ0iS6iIQuKj
S/4oovz59STFAEyHDV2GSV7MP10wY/0L+VAqx2fRJzcWMD6ZJ1i9g6ETELjrDzrrzbT6a84SGuN3
X9f/AvmY7QwDIPJ2f9rz1R+8DM1Qw+MA87oeWhFI/fgiyfcgiH8iQOrRpeOqJowEACxxQCfXGt8/
ZPy+kN01uUobDFUq82vu8b1QCF78I6yKqlVr8Fc5xoSpXscqNGrCy/f+4uYghmxnsh2imZ11NYGW
FEDjSGtKCC6ozfWRxqVUMg7cNFvvoONCJ4c9CHsBO8X5XJrHVjO2+YrCartegsqn81cMyj73jqJa
sc3+uLb/ByWxAdVvIVJeaRlyaxUPHyyWOUf6E9ApdDUpniu78JugWgMi4huGNFJ9TaH38Bup0aDl
hxfX04sSHHHwaL5I4N49t8RJhpnbXN6XXe8Muwa6LLb4qhtu1/FwfzvnOez/sXOS/I2JCRfrgeOs
SYNZzUglfrib2k1Cv20tHZwVxUQa6PojRpiTF4LIc/hCBH2thNvXvzXy98taY1VaxTHYllDhRpsE
OVzRmYvopcT0hFGgTza/hwENJEAXheOMm9nBhJEwvQsN9FrKhgSOXqEDBCtbarSl85jKrzCPayEU
MWJojKLVKRaP+lnY50aFXMSsAJhueddMaKOOMByDpqUp7VYwr6FRg7AUoLMoCnd4ecEYDT09wnGW
R/+OvBJHSktxVOcAlyLW14p9ST3mB6GUEej7ZTs3RLRYdav5V4cQAeEXmykfNR9uLXY2xCGqwut5
5iHlQ07Du/BaV51fZ5PHnOH/L8iOslOtxIV9ShtTyXQmdUlmU3IC/bEcu1Jhnr3Sr6cc6GQTYMFY
ai+XFXtus9I7Rb2yWjeyH6QxgfjAkRx+3IMNBNFzLhgA9BvM0lDVCCNhA7f6NngDltgS/Acs4O4B
u8gCgY6iNxaSf8+kgMaLxEb0duopNjU9UG+Jv7UoYue9euKmioSamShBwlJ6pFplR4Tn/O5ZxO5o
L6z52EH+ErUyujEFXBn89eNZvQB20x5nCipxToSvdcuZul9BVjagaRyz/H/k+aCiV3JCz2PrhyLi
4dhagzk3iYF1EsEeKwFO6IPxzWVd//EBSeOkbsAEKgF5y87i24eZoSdu4sj7L5aulLYQODUlxHeR
5DCHWVtp/+sIRs0lB8IJF2+IGJ9O4+USq7txREC8kIqj7Exwj9E5Er5Lq9fI7fHxYvSebCObn4sS
VrXWlG97nXFCnTGazqqmTFitJHnx9HaboJUmORCvmmelYzk6+CpswxJkwrDniNU30HmJKMYlJgLk
KFpqNadwH1cUn6EE9z800BKY/W4aSnY/EOiTk1tHs5aJfejV7v3z1BWZa6rRI1hejk/cQtLa1xS2
cKNcTTpr8P2pSFYToxPsaHtjY/PrZ3XNNpjNmZQ0LTXzhMc8TaILMo4nRgfyw8b0IjwNrxD/wybd
KRVieKalEOL0EMB3gvESPvXEjjrwjamLVvN3xs5Ajeagd5llDlg6S1PJTEY8xNKcGd6DC/0u5FE7
gqLlxlDsk/tGdmx5ShuApLQ0rWoJP6ECatTAkhEFiT3kkh+DPEEPUrkFU6BwHFif9yTWXkUGeNAC
H7ve1wGr5QtvtT9H3eeEDGdzGuBXxb8lNRJhtOEyB4Fph4rbba1Yw1RbjtIKd0PXK6LUZC6xTmq/
C66yWCeBi3P6+pr5cpeNQrfL+7EeXF3nCNlTPNRTUJN28iGgt9SeE3oMg3SEac9e0mPwjh5uJ/4b
Eug+PM+lL6XpCWoCWJ7Uw8lxDnPQDJf34UHe7eLdtRCYJxCdIBWL8L5qxzRJPjB3wUL+sSg2fedo
Z5y3Kr2ptamSAFKr66dBmME22ZutBvL8W0xkXDbVOufWfV880h0K/xmL/yLiyaP7uuR7QbEDdcmr
daM8tI+pgN49VO+z4bZpX00izjfMAWmk5VfFH492+3xuAOihZYxm3b3a5iYZ/IsTm4nsHPkMSUcV
Wlr7/qf2hOImjQ9rd8Sra6/EIIHg7TsA5lC7LmCIUj3Vbu0KZZxQ8kgnhc8z5VFdAAqcOsetcH8V
n8y65X3thOh7PmO+nkRtp3BJj8yfkHoTq+4oMgjnLDvZmzOVsvyrsYwtuvCV/qdXlabqxqakBbQ1
4CQP8l+adhSdwtOXINPDikbn3mCWgs2F397aKt+i9po9X0B67XXJCGrsicXJIe4Y8CXTTejLwPdb
2vOGQO2gjdikuU1ux+HbYLUESgezAR0ohMx/U7nafNr8+AqFlDoBjUJcno/ZWVzrKyX6Al3urNQS
gTkRZN6p+1re9Av08oUFHs/LU7J8o8O+86xRX3oNDcxS4w6vsUnIzf0qZ+/2rCCu2At7389Wa+xp
mCHZgi3PPCWm0gJPBXepuk/4eM0AEcyc2DSaMdOYUOz+PTm63iHVdB2qt/inRMHnhhViKGJk3fM8
g/fUs06rdGv6LyJ4aZ8iQqyQPygmIeoKx/BEZ4fRgQUqesREWK/elj9f+8thAPlMGksqlCDclznC
qwLy9eLsCSHGEbF1KfjfyBbg2xvg217ExqV121TmD/064bWA2C3Arxg7nQIGsEGlaq5PAiwcoyqg
3RgGbkoxWMBq6wzC8caQ4YmWX3FaqaVHmzKr4UdrBWFekjxnyCL/+8jXE2quNDacpuf1UKPgKw3Q
40j4LF3axgEsrD10Wx7z+vs05kdloc30QbU+BGeExtfhXJRY7B2GS795ou9MJo9hq407tjX930NJ
RWptVK8+nTA9IFeQ2ya58zuBCIcCe7tDlACIdgV3X5qIsK8GoRW4qXT+eDA76xM/5ZlqExnzcRPe
aNooBWrCo0LJVW8Zq2y44oNHe7inA8k/Z4pUbG+vUzIFu84qb8czvFw/EZEX5yOSsVjN1UJom0JF
kTvfYvxKCj54oy3WWLXWtMMJ4S9SffvhUn3qVfQm0cyWlsTs3uHdEue170CsGJjA5lHjCMpNvEmn
koifmQ7tk0NsUwVw9AzqNDnYGJCSMLaGjcogFuvLw316o14b/Vfq1L5qJvb+8qRP6n5hHhzpVHHs
K4XL9h32e9kop8/KqgRpHL6m8c/z3gRT02B83nEkqtrvnPlg8V3sPOo8yhjByb1LrqjTb536PVM9
QDu7HrWnQinJoPwg2ZlVcFcXLamMx9+lG98W20cQgvs2PH4iD2gw64zH7qOSulPiIAWOd9GVY/nK
KCKgNGKaB7J+Wkgnjg1esa47khxe9XvMoAJfaCMDtErwsWubfAfSt5LbgumyVn95/5FOWRI4oCxF
La9J9y2Pn3B9qzWaZa3Ete1a0JSyVooxtegD6pG3lia/6MVP7ZtsjYovviOg4dD6ybUVgq0HPjSJ
bD8vyEAcuBX3JkKAQPkLH1Ep/ot/wlSyUSVrrjfdRaTvYfp0id8Ea+yK5lVk3+j9lGxRXrCKuRtF
ratbw34otTKrjjGuo+KQ9LDZeW3lytvBirhkfH/1zfUkJkCoTS83f4MSrnYIotaZ7ON0W7iisuk4
7Lwh0CSNqDPcnxAD8bNVKO/j0mtNtJWvlnrKtcZTWrOqeyIasPokurhu4Cmymo2vui+8wcSNOpqg
v8d/UIaMJDRmuAC14GV8xagRmbaNSqmpu88WixmVXMciqhyXAzRsX9tZDSUa8/nEZfhmBnyzVccf
tUV+a07rUR0ulQLTa+pj01D00YkpiWYR2iFEwWkGUqV8yY9AhU/6pWk0ZlsIWT3WpTu37ZFOK3o+
cU5zLQDgKwBwmTwaW3Rs8/IuwsrrCbAQholrGyD236ieDvg0a9qfQUIYoLU6CUwCV3aF86Dy1N8F
5A5Z06NcQUD8BLqbe+dPprFInYoScdcHWH4XZ1CvUydOIGlHRJBUGkJi7JGEnotehdmgffwoIfCD
79tPUOc40PGioGYGdWqc/qbZvF5y0Bys9hDQ2/5y1i3KYFk/3Uid6yycdqNtCP6py5y8RXWX7HHk
FUA/Y01py2U29F/hKN/idWDfZKqPw9sBdSQ6WsRZpZWPn/1/SN3Xd2aY/N78TvUaE26Zurwwy602
HUQM5kw7L9al6/+PCn9guf+1/hTnerWYPmJkTeDLll6AaQXeVYv4F8NHsfO2uPk0ZoZ+v8x2Cpyt
mBHPyfJcYeDJvg3wca0Laa8RQk3JcPxaCSB8zk9mNcz8fYNrebtAJ/SkD4OtqEiteMMJL5r/igEA
rzb+XchpaAfQHYSALFk/GpGcQ7AiyLHuXZKnUvWixgoTF9Ayf3HtiGzM/Mp+cOdcjyXUBDEgvf7X
qlk+jL9Uys3aC7wwTiTBSWKuknvtbNJESAzgDjkHw1ujg4qmKd5SUAWBXmKmlKco4Lz8yAu+J6gw
8Xw1IZOUPjAGtVxqm6KMDYxG9S7Bpiee1SPx6hYEgLVvRDSoAlxUjpg0P+L+T96wgUniB6Tml5Qu
5r8c0Hc2uGV2ug/qacWQuS9ZvpLn3boWnfgyjd2y8JEm92gQVoauGoVILuKQv45WIVxCsTJJSQ20
IzGe1av9BrI1aEhbNJF+7y0fIp4eXTa62tTYxupJDtrEQvO+TAQJFaNekFuGJ78lEYYaZu+sWbMJ
MEoC33kyU/wgCAQVgDFFDyMqod1vmCmK1ZW4omdNLsL7yFnT78Bh9iylwIOxamfPwOXMK4aOI02A
im5cWI1aEuRdja18jDa3g5r3af6KlDjRob0SFGMHMv0xzT9S5+QuZnkCTLycB5J5EHlRN9OyBcSt
qU4VlV//FW3RZH4LlTZVc/5o9NExJPy3rI7SfKBSXmEYO30JYvzpXnkZKK0pr6AQo5aksnU3uHK5
SKiHDphFZUQodQzkF7wv+OoS+dAgJuQDs9YX5CyCtGGP9J2Rawj0S8Iwqth81z/byhb//KHNLjwa
fiti4BinkmKrg7+Wa9sof1eHAzAalBnOdmGv0gFTE3G04m8dTn+dmmqaLqwnSqtrfpwt60JOy8Oo
HQQD+Orepe2o2gdlvR/jKmOQrjwdgL7fGlGuYF9jVuNZeWz7qTLhwcrFM4DKnhofGZsDxZIJamdv
bHnfCy89xzNUyGuM0c5nIX/zPVNMk2iIkv3KnyOIDo1AmHn2xX1sc7vR4Zv7GS1skTrkyZmYkd1j
KtxdEWP3HAkHDZcCMgKCb5z4vSjZCDMQn7V0tsT2XoalagPCmKF8d0U4zDz1MZEuYwbAIdMsoeNa
awuxTJev2dWfV6SYuFlVEsqM55FM7YqdQ27tZjvZ7lR7vkTocgFMbt14tpyCSlvyXcQw8TloDn+/
ucH5xbSTMkzFQBWvPE5amo7wgKHuT4vI0uryipu5l99kVwlnMDoRjKnXBOHEDXZ0N54y098ssB1x
7UJMaSGX13Xwl9RoM+v3KUbnf4gQFr2PWzD3nGSxo0T8oxWKAN72c4+chaIWIsVsTV+EusFjmJsv
AcWtL73cM33DEaRdL8rwCp8sCaRW/QqvAb6uwoaaFDB2NNz1Hxc6t0uX6silGgO07f/cW5yF1bee
mULwrHLhIaXxZurig0qSl7DYbcXi4T2WyoAbFKdIOL4DOgUyFt8eIO+YDF74mjRZRBFU0I4Uw6am
6m3SFiXdF4YeVBuVFVyZds36lh3Soq1LkraS0byGmSycQjTpFxeK4JcSvIzR7M/6seZytoFuMbLC
cqscQTCFQXYctv+yLqgdsw6fR5pFElTHx54pBGoJf5w3qwCYAHd9Mtj04+ZCafibsBxzqDBBTvZB
X5coIYVnzuwI43kkPr/RClKkl53Y0sZecf1bdAHrelvkbQYzRWailUt0t/z6Xe7X1U0D8LkZ6Cxw
Ep9yynQRjnvAQ3RM6wg0tvWPESjvSpEYnRgkvJCseGW6M0O4VUdGQu0wS/V7reNuVtRB5iRn507d
qEb1svVClABStiivnJD5n+fzMtf6h4Lk9wvtZj9H6lxGnVvSu2xLbQKkw9YWqz+84slQykHGoU6u
SPw08K0Xn1kg1bRBUlpOZ/FNzXaSC29e4eM9fxAokBhvr7UQsYv4lB6VFat0QP5aX7CpOfAb3FHI
OMh7LIUKaeinx5Ew4q3iXqZfQHGYVljk+9LiaG6dEBMjz4sBgI49/SPfGJwaR1ZtMGSY/k+FgJYB
6Qn4TeiyDSdEBj2tkqSVMVIoVtITFI29Y7IB89968heK8UC3w+XdmAPift990KoR9gMxRYgL6m8D
ki+dGS2PXPNMI9ex+6HQN6IjoHrD+pTemUMSxULFh4Vf3ffUwB97XbDq/dRb78qaBOLn2EwCX8LS
A8Vul4h9IVyONJfbkMjCKzDM+To4F9EAU2mz9BKDDPD0GxyrfnMDQMSQ8wXuStbItt1ejTMMVmE1
K1L8zxU6Dz9wBT5GlcB2AxQWja3kGlSmsL9X9UtE8RyLHOIPv+AiMWzObm/mbjIz2YTZdT1DjSp5
bU4TFKTDOXLfcCa6nXjHtLop7Gas7NHB4Y+IDrTi25blKwFqI7+f5jyB/gklA1iOw570VgS17gxQ
1sP13FPACxhl8OASZtyBarQIVwfVYfyC1lN7ygY6PnSQU5rxBQeETUGl7HI2+2/i4RA7v80KCP1x
v3T1+/RK6zHAazDXv9qQkUQUJ7DX3JuLERF3hE42x4QImWkOcaKHNsRRLD5TJmdpkmIObwvrkuq/
wu1Z/yx4NY/gCavFNro18XENSZqX6CtM0k+3jTIr+bAmzCs0G/sqwolmQlZE7iPyxy0xsF6v2RWK
WwDGqZ89/IG4B8coVO3M3xhcnmqx9/0n0/IBdQVB/qlDn8dkAcbTeWv8XlKCGE/i+tZcjtVkT7t8
RuPZjyRQeAj7ieQKDwMa7myCCtzkTKb6ig56CXOP0xHmT9FhPUqZwVLn1DpvMF2+Yw9GphPpvztO
kJshi6RoYt9O3RyqPgzsUmcm7Q1mFP7gZWrxujKZmvbtkBGdguHRTbzGy8tyOM1/TL2ECFfCeL9N
RKlB54yFPmI5FVV/2ib9AkLWAYKvOD6z6JsVB7Zp1MVcr2Ka6MhkGsE4BR0dQaTwcb/vKaGjNFpF
rIwnN704/DbSKXQBEW6AprCJn0SN0IOFFiN1Pak9DMPKQgeGQxSeZZXejqwGUJCYeGqq2x5Og9ou
QFov5L7Y/z8OSvx1ule4oU3E9KMPxOSpPXDnml//TpscQ/4g+p3jFexclo+Sc15+OvzV1Etya3TQ
VU+TCBkYNHsIk7UUM2daczVBZFELtX2LyNAiCjTc7uPVsHo0AcFVHRK06wZF+03MZT6BPVNQjuF1
wlO5fSuRG+Kf6Qoi3EWF/B0JVyxQUiKPR147i6BIcjaDSchKdynZHUi6AK0yZlUX35pMTFlWustj
3fG01x/OIYbsXrqw3rQdOEHck1sbOsH1w9yEItueGB7VVrjH96qxXDtUBSKge6hb7tm7rKR380Mb
nQkcH9yFrRANf/7wlSouo7LypiCTC0mVyjlYeAt4A91UXuUZTnW5HfaeFsxO+UeR+Pb8dbVlUbjr
z3iRlqwckE+kvXDe+OkuKixcEV1ri9PtxqWJ7FAP3jIsUZCxH2y2FFM+b+bMc5CWUigYWNEntxp9
1EdCCT6NTGsVzo50Ja8kKWZjmaeE58HYKcO4LEpi1/2BK9eSLYkIYZikpOf3SvVHb+H2uMR23dx6
Y+EgBHz4Ch6a6B6ebkmlcgo6yssTzaHXWs2g8u4pK+T3OjxM62w3iJ+Qo+QAM6xwM2Te1xrkADSm
RxLee7tvFkUrV8X24ZiMIKG33xlzys+ELeT0RW3qG8+Aum/FepQ9qdl8ot3oGW3GcSDnMVFOUVPZ
8yYir8LDQJ/nSPwZQjTmHCJeWxLeq5cvf6ppqINLon5edEtbQn7ODBk83g4SDx7qgzJufw/5ni/r
bkv2LZGaQk5QjserX3s2Rqcqevdxnxb3VNBCe/LXtHMdqLpeO5rfxJMNaIgX3xlD+r5eTSVEcmLc
oefjVPmNOB0Emjo1A4tk6jCOU3M+7yMbx2DFLpSUBq28hkH2zwkLqkv6wQQZDBbJPWpHtSTidUID
dYEPAH6idFjipXSYPdQuXqfHhtDVt+LprSiAqcQ8THM/Wj8Yirq7+APnoEEnMvmwkXjOfQLlIkoU
Zq2ncZW9IZpQyitJ6VBn3Ixzk+fsxdZSa1GJhvzn/3fU/RKf6JXPlQW73AZPJWEBuYQacRrCTE6s
gkDBjtmdQSebAv59hI9uxihMIqa7v22jE4IEiTw9nVL6tu+n2unT1tFQSFli7z39C8mZmJpI2nga
FBz8WmK1k4iovtDTu0DhVStIBGnto7Ck8ZiA5pB99GMNjNLyihq9nYzEz1yTL5Fk1nDvdRLbzgFG
x8/1C2RK1Xc1BbRgojlU+HVuOxmfBSVwQHbgMVrhAQMIbCkrppHKtefKygafmHqs5BRUh+Ee/5jo
anXT5lPzUoY9xLtN1bM+WVCMZnguwlW5sO7YNYKJGh1f2O1eLgDrZTehw7yh77Z1hGf9Xr6pyNGP
tqOrCJLxPLTCGCZCcIu6M+jkvcFiDO8tooDq15zhIDRLbccSIU+a5U85URoAMYlkBWtCqzW0UPWk
SGdyw+zgOnWbTbZGj/79YwCvbtnC6+bc4I4Wxf3bcns1tPHpmYnzsGJuQITK84Wqe6OyPa1wf0b3
y+an9OFyJuWAyUdXx6RXhKnODZ71mQHBPnrhgRO/vVBpNw0b8gghAhv9f8Lm4x0ezvQnGunIaCg2
5vpK6PhEQMcyaVvqB+UdSe7x+AGJJYdMaknUio4JIxthP++BSPABSZOw0mrbd+hVi//wzwDBVlZT
sx2aoArGMJFrDodfn+yPhj/fnyri23GbFA1jR6GUaMWTFDYQBsNilIGLWeqSaHusRkTtOOJ2HZ9c
vus0MOsWUSAQmwJskeRRbyOZA3Q0I9Yys3oytQvqXfg9k5+cVCwFp0oB773DKQ+thkxcOiLQpKCG
VB+n4bdkHL9pcD+9iavJKR4ida0hZYjiRi4+O/b7eNn0v/HESf4KlGilG5hpww8+tQlDUB8uRGbS
gSUPkneHELxbizTkIwN2WWNvgnGYVX59E6ilPP/OZh8AHoxdVMaANZLFPf3+kdrcNfRTBCmZYSZ4
0XiV/L3UGsuZkB1KmWyz2q7g+Ts2edUjyN75AGmLE6pXylxSCGmAncjwgfptY/zWXALhXsIV7+cw
bGWBq2FJH6fnV93zbZZjymh55W1j78MIuhnmDT51JZSAyyLFE1sGJ0ujeePYykQbYTUpXHXwbj6B
NXwpa1l0pvP0CEoCoP2iJLsXQpOgKMiCAIQL2yJEDWc6kPz/swCliKXs/o+hYFfk6o3OTeEjgj4J
xdzauelEr/SJdB3q+Al9j9OWbGYXUbqWtoJ/4TSX/yJTtoIJPO/8XVu+FpZgA6ZV8x4zFOV/LDpc
DhuBt3BFOm4aAOIAqRp6FkXsIN2K8idoilTlopSryHcxKGPOZ2yQuwI6di+tLnNNz6pkkc4UCt2S
CY6BqzKcj3LZIn3hWTEEn9GoXc405ChBTFckEpdR9SwCMrXc2yiA7Si66GDabEjYgOyQRIZ3FEB5
8AQh6GPGYhbay7pBdctxmO1rLmqcPo+a9gHoUZUP5efSimtuZU/OgsHY7unNMePT78yXYHUb/ME/
QRSsQZ8tkmgtUEpNNbHk6M7miJHdbM9tGyopOxhfZRxN4y65N2WJeJ5gGyhEOInJNtFnidBhKoWK
NAmtV/uvz/dkjG6bi12rxv3SmRXo31Vmi5NsXi6FfqTi6+5XhmFWIJc/FIMdr5KJYI+XWpNXC8dy
C2Tnhds4rbwDx+2+9bHNuEuo5YMG2XXxOqvVPSx+N0UbcFMe1p61kph5J1Xj7tVTXjUxaSmWmLS4
Sk82m1HJpvOhV69Dlr8UPRtIcPfOyd7b59oKZGC3t5g10WYdGDVZXE/YKvXltSQ1tiS/dpwNzMF+
SMvjwzOa4kzjTJ/RKoU2xe4KnkSr75aSmJMgJEEaw2a5TILXwVxwAljV6cUU15R46koEzHTaHJKq
Yl8I9nsWugGWVbbzQP1hPEu7PwuTU4PQfhGXtSpFyb9uJg3MfTkJ5wcIAxkXkklQgR1PepZzjzbb
QwXkp1P2EkNd3BIcn9gCi2Fmuv8TZ6iCpkj2ZCxZdWACDlNNgHsAVW33PdRohLnIwvXvEFernOrQ
lHhbboQ/0VufqXc0THBJtVLSRhiVGHPfu/fsdnlXBEsDYYGvelVfugQoO1CXwn1Qw5NvvGxjpnMX
P5Znuajb60YRsI0k6bhCgF+maB+AByEqyW1d5araXiemvRYTIJUfbV5XGxeUY4C6/JJ6ZrE40C/C
oXCtyrfBVMKTomLo1adVHZ464yJuY73AIsYnx53OFlQin82mfheamskr6DMeQP+b8SmSn7Lsp6z0
WHHDuJgBc/iDseo3wFqtrQAvzP4AlcDgfEJzaHX0S4G7SFdk8ci8aAxlvhlc/cClYOq1GBRVS0Dm
M2GAeeirijVszK44q49xITOHX9DIgEjg6z80eP6hPvmTn8toNmjVOtBQOO7di4DquBNTTYtVEdbA
8wRUKYfbVXVRgKZ5HB3YspjQAlDiC1KqdaQHFk6c5DNadCLI6wC2IHCIKSJpcwM6HzhS0KWmUc+H
umZlokwkottn0qz0yktG5vufX/QCw3Bau/p6CmziEUVIHGKgNHxLSc29Zp22qMnEvVLzNru7qVQi
jiPTdXjzSi8A2Eyq2e4Tz71dkK8NLGNV32bSNfLxTqOB4bXx9tlFPJ7PpOOcztx0mPCRF7xySNxS
SA1zj7y/Kz+it0+oc2riIHYoYK+nGTGbiQPv91fymqoKqw4sZkk+zLduaqIFP1caWCad9j7pY4kp
3B5fv9+8VtkXu3Hpn1Y/cAKD8CicYeTsIuTUSpIv63jhRYG7bDKQoJiXlk9s86M/AqZ/u6FFK8rE
yLaDc5dPupjtOYUy4PZeZdgyJzHhEev0wnjLOBuV/aFxjAJlMEB4hEkyhP/LTjACVL6k/BCWMiNT
fjOGN1LY3WoCk/moJ/+Q3B11aO/50XDBP3djo9oVil0Ie7DvbxQLhZKG9yx1vvTWgzj3NEOUCkRY
XY/9wFy7W52QfiEfBtDKvRtftkasjFvAmt1Sp3qdBVLlkaCqzCk/o9qoIe1PYdcfUBKfB1geGgmk
pd7XdW7TmDT86Zsl63zkKYT7+AEMEj90sVvIGELnZ6ISyDmFNQfnF/xNo7n7/OI3PzcLgg2gzaPe
G6rUVok5eou5iGgc/BxqNG4oZZHM+fW0r4r/87spfhjZGtU4EEb53oZvU6nf19tiM/xMF3xaAEDB
AIrg5kF3xSDxcsicgzmN8R0jTxT0UuKt/rDskUj41boD4b5rROwBO/jBwAsLQBCQp+sIsfCEAnq5
fW0TMSksVMSGn9s19KaMfybjuGhXcsVwq8VKK5MmHukbexFoIkID4ZWuUoy3UvsG1aueZo+puU4T
b1eZyJlsLmtdlNIKDGRLeJojTsNqK+9QVp7KdpzGDkgMSVww7qMbojZQPNS/PWnNUjo4oVF4MknO
9/0qICT55BAYF3gA2Lql1+Q+/+7f/47hfSTr2ZKG/4BONMzvrf95s9ejXN8WiYvEsUH91lXWl5o1
CzARSGQnaE7rHArt9sQvp6PBCn3kTZEXAlU//D1ln5HHsEXkN5pyAPvMPyZtqTyfflfIrMBHCOOr
/SCqhQgDaHg/FBSPkeL27mmFkIFX89Qppo8IQZWpn+opPiK7mJoIJj2igSon8ubbiyLp9zrOGRME
0aoTDs/vdEBILttMm5834mB0HDhLB5Ek+S9V2jow7LzUxE+UyZAJLkYNQtevflEyvMu8agqPMPCg
t3yyrnspKox93V0eH1N6M+BtfPDO/49kQkhTbCw3rjcLia4ys5/ckwJopbfume9win4Lx7ZE/J2X
TsbNxkNB2J9h/vIo7RrAfa+hhj98FlPwGMP5a/LswaAv9o8lTpEH7vnxu5mo5MFHtVWOmjNocQX8
kpz5yQO9kbFF/pyn8v6JJLwkXqOYlMvN58iZ1bhV6EQ9WYVNNuOd0H9c0tBoVpmCUluok/b0Qgd5
UflVriYUNOz5twybNNGNGX5fppXf1BXh4yx60yykf8/0ePKSkpk/zOCSigsv4azSXA0d1j3m9DWw
/+nqjgGO9gI1wvH3PjiQKegsLSIo4WQKuQqvkKpebCC7vgTKXdHZLp1ZnDoqeZ/NwOepU0dSycyC
1Sk8+kOqN1TE5QPSi8EvWkcHYrlL79K27J1/6nK6/NS1lIuWhPQgyvomDTgq59R771yIgcYvV7eL
3ACVM6TgYXIuC+VUoonYLxVdnc80KDJ9Sq2VDgs0lCKnyQfGB4Cp2wBCJt3WPrHWFDLU6s7kw2jI
6NaooOLKd8sWgeMqiK+jNlAKcKUZhZtYNo3SzdMOoVHzKp04pK57Z+CaMvHwuNDbHrwg8HMo0oai
5ftiPZnq/EVQnrAsJFY0Vh8AYQFy0J0BotnR49tRyoH5mT31ZmRWPGVlnztMLk2JK6tt0UjzYHgB
Od80Fry8jZf6LiNkVAt68cZ345wl/XwBcOuNTqaZhcr6Ckk2RBsviICWPCuLspYqT5RXTU2Cr1pe
1BS2MHyz9PcXFotI72FLiz3eLGvmlv3KTBcQpTTGGLqwRz/lic2++FXxFnmeOAq9e014MuuCFfcd
RqSf53mXgSMIQsfVf1U6FWW5TtgBjzKEfb7xxYFB6vIMp4E1ghEMdvT6WWZ8lRuUsuE05jNyrbpZ
EpNQnsorRUpCFv0DpYOZwdOM8/pV01WTnyCQDcMZMJyQBPwo/78kfARJPGfK0XU92EFBA8g0vD6/
00f0eFEPPF7pdaA24IwwP0WSeQSYvsk5EdNVj38uhoMnrsI8Uf9DGqYScNW4rrtBVdG4vVWIt+8/
qg1LoojNh4XtaYIE+Ab4Xo/rhtoEjkzpCkqgoWCyWsQwYpfJJXSfWXf3uVDnfuLVL7Ik2Ij+S0mh
8gkTOFIU1SJaRIgwUkZ/1PDPNCsdDue90hoZHODedum3dEWpHCqh8Yar1QOH5GT3THZHtpV4CADI
LjZqHSWT4SOaTXiH0/tPjG47mYp61DN1W7m7flCOG1EZKRndEuNFPUOLCUseVSVjpDe1wbpzrH9q
Cv9C1tYGAahKbNB6D9ihScpik42IAYF9ES7//WyhcW673gd9sT8jnkfTbUDXD8m/YWYKs/yAmvgk
Rvt7D3YCB+VDjWIB8zlco/XN7w1Pcg6uaRH2P6iv03MxtgdWMIVrcv5FZP1gdfcnHLZTp7O74riY
QWgmlIvldq1HZwBjFsbfMRXdbIXUFNvIRgMdePv4eg7oT10QG7N4js+ab/hKxnWzVF9A+ixofyMU
jEpPdoCHFKww0n7tXsGl0fvOAfnfWxVtPYvd8cDnm91wZMCrzvRt+7Eje5kXX3QeTYcryH+k+hA2
gq7GQo3H5yxEzN+YbnQ4DDO3I6iamfHB6dxE8+6xfy3l+0/bJhnHFd8HJ5lktqm5C06hURN9IqWI
ovQftxXgDtQIP7Iga9KmN315o0sgBEj1RF89+kFI2fWeL+akxPvVpNKhL2QkLavCY32siXK+mdF2
tdG5Wv9KnTkp344mGeX62ZnAgoayQDQu3PeU5cLuu1jAl3gABbNvFFVYCHmNTbdzKqqeg3s2OfGl
jJKLQRpKJ6tnMPXGYFXPRSaAm1MRDNISJGjeZrthID7p+a5rP+dBKPdN+AdfbW2YPx/IHR7BZsLc
ayXAN0Kpp5ueNnTa//V0X8sAGuENGe49XvMDx8Kc2E2XP9pG0DUFxqlY+sWeMwjdDZoICRj0Akie
Gws6GR7KNx5yu5JXBTeplESfd1KqQrRj8wh8YAL20Qtf2Gq4UFEf+Z6IG67mq4b2UjZzpljj4H+r
rXo/CJA0lUcVSJmCpB1WSIVfd6T3H9nN0X/ecafEuxjhJLn3FQWeio8X7iiHwaWk1/88s66H3RTW
D6lEB6Hi+gAEJZDThVn1hBkWfpuOS+rFg+C0PKb2VLqLxkH5SruZa2LMObBpSJYHBMnrQmm1qrcE
OXxeff35Mct4dXZ5AY1pIr3FpNHMceUAkEhSs0OV8ciR06jRVXhGFIy0P7SEy0AJBpZpeMC87TcE
VNmirTuDREz1JskwoekpYF0OkQVXXTxm2WcOoNFzcponCcsE0XtesKtLg1xkqeAuH69Rk6YSwVBq
HG8fzunxY0ClPV8+Qr3w5uJTuUusBIh9VxNTblrC5K+OapywBHu5dOq+H4DPOGIv0IHF4expHdNz
NoAr+jv4BLevV9/jn3XVDhZMQUeQ6V+C1ktW/2ZgF9vEbPpOap/WQGGguD9uvwSryUiOELRTA7uC
sy11WwPHgoGeyMH+Lh21f1VRuDTnc1dIwtdyoaQatDu3/REA/ABDU+WrftzL58Lpm6Aqe8oXERGC
LoYFCEFoxwHW7jACuD14wUKUGg3RHcGocHbp0o8WfvrUbTEo80HX9Q9ECbpov3/mEEdZ4lpIPAH5
Lw9e+zn47+R9KH/RrT9iRK8Hi6UTZnW8F+Hb3EKuFenxa+k/ATgPNC5bxtUq548QbwT8esdcsyAj
8kHtbdklyHAvGywaHqwUsKJUdfxWZrt6gRv3j5N5NHt+i907ChM5IST+V5f7XFPWwleEnYglL+MX
thuPTWT5mgW31XjXk1x7xgv0Q6+07Bv52WdNKI5z/D8g7BLln5EI/XT+OSmCBrlSIy9aNlE0q4GS
PNjwHDlB99c2DUFhbDMGwPB//Ex+6Bc+eX5Y7PTJs4Qrma2eZGPt2XCVqFf1u5FsCggK61kXczQD
DywfgE9vZ0i8iUgukD6RKYRUviUesT+0nR9vxCqS95LO5qXTBrMFxM9Yl0OJv3pElzoeJ8rX8CQn
Y+r/54x7uSopyrHZ+CNIzCEgGctGZu6VsKa6lF/kXCtOJBBItsJQu8Ew0Yke/yq1aHgBXW4Mc3N7
bR31j0YKFFUsRESUqzCbBUmvTRMB54VgBarGADebKrisvzoTEDTmvRo0CiZjIKn5zN3PqLtMuBig
xRth7efp1ba39+qCIYLHouuhlzYPQmvLA06/bwgx5uII3jeKLAM8ZiyUuubjXIo56FMrcK24fm+6
t5XRHlWl5T8nVJQNS4zHJPO0FwcnPbPu+Zc4oW8VVtd5RSy0Cp2oxsiVRufuHwx8t4Px0x7Gugfn
1AKBFGaOKENSJK9SOJpVqOp+3E2u6I5bSwsEQNaW5J+JkDwCKCz3VOVzrj47n/OWkitwpMKJPXeQ
CDpY8DJg1MtBKTDP4qB82Nn3WiavzFz22kpKbAE+hN5DJwRQUwiC0RWbVdj0OqnIbWGX0bDYOmZG
XySC4ImWQMG3EpEMHIbgiwnv+GblymPUc4LmEUKhhFRdravTUVhOhQLKRwTGxPTtFSD98/8yiqnj
ZQG88rtj76h7jArg6aZQV7+dCBtnPQ5Tj9kDXgN409pv6c1rFViUSPOiJWai1aJsO6zURjW9QsQ7
jPQVx3N9VFYbTa/h0mdJkQrD8cw0mRRr1PjuUGANiKM1yPJSk0JXDYnBQC/N5042ErKhIk61PigN
ppO0ycEI/Tj3nC5L+xrTcsigsc8R6dHg8UW0i8c+J2FVGWxOthkScbAG/gXd6mLfyjnTo4LoRStf
l+ugC7FtmaxuixGSGm7giiWXtRfkt+pC1zeb/MNPOJmAzebaNgif3xqkCmj2b94Zz5DPELaHbBTm
FLqStQ4GXZ+whT/QiBWYlU4hPF/Nz3+IXU7os50LEEFNBuRVQztBKlHMDxStwpSXpek3etwF+yy8
1buwwu84EOZ6Y1RhxaivYiRESDx4svKc6o3tKVTFRCZiJilI+kqAFluwrTwR6JNum30wnoHuhAOG
eBRefP3cY+0oHTo0lQsq7+r4ryZmiqPpnhATaHMmHeh3SKi3uaHnwkI7FR0pXc109PVKpiqLjKR9
0F8H6d6b56arU3eI8XZ1aO9QSi/oYoISheZmtVekZcBlZN8QvMPABbrjLiFiVMvA0PyTeyojPfl+
u9DoPqd+DUb8+fOlvqi6jA09EbJ31XS0TbuTvUIePL6OXa3Ff1Q9XteIuCgefuL7Z0FKYgGRP3vo
sECFys6CggRTpuIv1J/pT9NAvFkaAoIv9lxv6K6ocYEP8700QRrUrjrtIc1XV+hc3Wst5ejfDKxM
fJeEn23PQfTC0Qi3qrbFC0zKw2LXuXJxhK1pTB/J1FDDpH2rPT4P9k2OGSPPvFiy1kT7StgdWWjj
WBUuvyrB+exKWjT/vv4CUhlHMeISh4eXY6P0dnmPxqQ5itg2KqFnaMUfDldtwdkQs3tu62UuL3H9
g8ULVnvytjGY9HUNsxWqmzu8c87L/rC62w77gu0lvDhwoftRseP8WUmPCqj6pFNsjTxMjBCTZdr8
49wHo22IX8QUA/cdO2zsTdYbpTu2EcCRxwU7X4Yh89nTfu014Ob+GV13O7rHoz985JFVvnJtycwG
BH4aZCIIiD1qv/nsZwCqZdPjkEpsucqvWhlzVADPQSOs81Wp60Pmh8YcYCopEjpNux2KxQwfEo/E
pFYmsH/r7tfG7iWyW66SeLr7q/eyWsFlf0GPpNNMcyKuBHjJZMN0VBF3sEbznsYYs4WpPm47jezj
Wa2wnTJ7nDhcO8ERXl26Q9Tg3+bwJm4MIugqnQg/2QRjfUJZ8lfj/juRv72GtAEIbsErsjdyChuZ
42aCp7TA2sPAh7VPMekkKNAGT8s2Aebvea1eBNX+HjwgBoNfT8aH9c7q9+B7USu8vwjKeYI0eVtP
9Rw5HtrjdBPYGD4W2mQAdYPNXcxRbV5+eU/B7ZboWW4MUcNEMmddULt4O1jBGVmZguN6oTB7rviJ
IVegLcQG3MWnYlNR3DLZq8oaw+9JvJbTrUeKAGcdmZxSzZDsc3sXcqaLHY+jWNWhVlXu3hV4NEEQ
hNTcQENMTY2GFs3PsvYF6+yD2tPP/yULPQNMR7vdzybR0slK+89z7FnKK07imEXiz5YKOabrxEJW
XQ5H/aXWsR7HKihcFeuvppADqT5Q0JH60LplV3L+zRuQrTYSRFVZJwqn6PkrTYaUXsYs4rdMHgsH
EtYP8DeWg7qOMniO4rC/v5hl/XgIHvoDdMOf4DYArkOUMo8EzoHEPc/RaKXr3DLTY80V3IKaaDBE
d/sl4Ck+5JgIe3HtA4DiqAtu9fosIikatSULMyp475mg5SYnZ7oYltf4gUGOlJOEdHM2YIQVBU0l
1LMbfmP9EOtiibCn6eEMSeX/wjB9Kr8BwMpCemcxF2ttTtEOqAEt7iVKgwYX9iiscoQNO0YC35vj
2/u6BqVqBkxXimC40Vu/IDz5hIuYoHnwPf9o10Wu+EMWSc17rb7zd5iEj+63xoqap0qig4hM0f5X
0Z9Q7ggxe2BnPqruVCw+Utl0ZN9KoGVhgYYf7G+dPya7mbOpwk1iy5DZ1WfOWPDDh8Z9OM3e3NDo
Ei5AmUoNLULTfimk4WeliQlvfAVov6DriPPWsKkj5gUvV696XKsLdHRSrnTWJelQODnsAfbw6mJb
vOOa/BULpWyIAM75TZ3tdz6uVWDnDGjyD5Ld/QQMhqK/vVO5Ym6DamSYzrB/31mFB/G+Q2FmOH9k
Hcl12Ili9YTtrwATJM1fipgKgNIbFsCVp8/0eGm039v+Ar+3dLAAjU9mRj2umhxlZH/llZ1pv6bE
/xj/R7aMhy3wlSYbBzxpLqTTKplS6YFEMG67QiZWkM73BoPblzom0N/M7jONslorm+Kdt+2adc1n
EVJyZxr9UnJykBB2qocotF2KUNH62mOjecFm7aDuKPEkHFW1Rm0e/elVLVX+ru6iT5Bc2Jn4XKcW
mceGpYbVEd8JaGtaQ57YUAw4RDwsXOw3RA3hWwNWmUqLVXRU68hR52W5P5qShQc1JfEWs0jFuogf
8P2JmQaKVtGc6fjJus8gTmU1/cFMnqFR28q3TEGPzxKPTOiqSmFnoy34yuXe7JYwsr4ieAU2zMP8
BsDK7fJthyl03l1tQoUPglxMl7T/v6fZseVsQfsKer/hM9T7FT/N0xZEcpk9kzipR5SlZLPizatl
ONyE2U05DSBAMvjqoGLX2YSXRUvl5ZHD/ZMBVwAWSEAY4vgne8Js5gJa30ND1Ni89NlLITm0LMT0
hLrguzgAwkn8jsWL/HGFEUHIbSiNHDg0ThAyi288vEg6qshjtsAS1J9hGqIxRC9uNAnlQYJ85ks4
0UKG+sBKT0cXQ7KBd4oUjmL4mWeoJ/Tqn7a4Q8SIXrpOb0PnWaRUsfXxRmp8dlY+jkAPz/O/xUkk
dV8YEZ0VkRFFhhypKKNZlkPw+qIKHbXr+BvaNHf/9PUjzuBbMJ63PmSggYowPgJd0Viv5c5Xy4G1
FNrGo5raHZNbQdPn/D2wizeWbbshqBBt/ELHAzipx86TE3svQYukVrUkTL8l+3kYV8BXAmsCHL72
42Rd68epgoXIHR8AD88flY39mUG9fw69RQtIqEeEL9IEDEs/UrfSpddY/4zwfjPGPA9yGdLOdJGc
s1ZfLtm9NjRODC2YsZlapPbZ3OT9Qifr8HhZK/GG5N6FgKSIxnrz8Wkx9chgeP1IwYubYizcT3Dx
lF+ZySYQLonZd6fUNxi3Ef0TAgC9Ld/1ez3O5srtzYwplT9qbX+dT/4IC3QcS3reTlmIbhRTuwVv
duFR7qvTx8+LpYzwkcTikOUfXJKCjMUXKeccaI08de2XRy2EEo0YE8TUQ6WkFmupCdVOj7C0qJmb
ncjMW4ISf2jtW+AH0obp6ADTAfXPqSMH/7KVX/0OtFEJSd6JyxO+qffEeJiq7weh1R3eiAT+DtRB
cEHolwxipqY1cDo9maSc4tBr8/XPU38bfUAuuWPOZAOxRReXr1NmPygRGoponztIMP37jGhP7qv2
/8qwIiMb9MRKs9J/NlqXnNKSgiAUs3z4xkzv+E+L7zTNvXbrHIKhJYm0+JwNVoVCxlYSRwMSS5B8
SIA427ZtYKudkDbmrNO5CgW4+yR78093n0V8xhRFMtJCOCDMWeQG2qPcUSshS7w8At6CTsXNkRtk
Th+eyLM8JZdWjksK23UwPk1wGXihyv3TVX5AkccHE+vyxi29SNFtVy4xktCounJv/nsdMvOFxx08
qf2XqOeDDuQwWx2fZgmmdNhn2G+8oCE+Q9EmwuiFs+c79/yFBqr3rfRZ+9eC0Ouyfn1vpcdfLDFT
nPKIVByT+cbNHKbujYVKH+BJxp/znRRdghIdPRS4l6jpnIP99hJEgckjoR3QqjSJQvLXJIydcoly
0BCXlapgWMq/z/acTyymcJ/yEuMnXOp65vzHTx/vdciyA6yOXsNvSit0iroTK97ZT2iJTMkXp5Ja
Swx2SzrgkBrAsNaM0RQ5wNxLPrcBJIJSf8SAVl0VooLT1OS7ZyvHihxZ6L/1eDmsmsAzpJUrhoAi
RI/awbLUI73Yhe6ytY2KxTpuckXJB4bFnkYk/C93ofsWk9uvKzZahpcW62eouPKSkFlWB+5TXQ+3
hsqIUMcLNk10x3c9UtpKTNCMAg5zbAIVrA4X/XsT4E2SU2URayj6kl9oxPYwdUvrKgPfYVIfqQnO
oSw/leZB4ABEzx4CjM1S/BBaPW1I/qqtS4A/1iAE2hkB/6A7vRkGbb8wZa7cf9vJ2c+JcZxx0EtL
FL4LfL0F4W5tL7PBlPYqQNCaD4Gl7NofAncHFFEmdh5KZKMsNv4S4yvf39NPV994fjUp6j6Nny23
/rFIsIvaPXM6SJ5MV4z8+g3JrKSt9xnBTj0N35ywjfMegoqvxaR73fWBJcC8qWhMLhm6K9x2uo7U
0KtGVM9b2Fhdsh4+nucNxdAF4YMOPu2a56mGbYrvtVTlJ+EeN2ZjOB/JSHci6dphZscm5qShO8TG
vvfmgF4WyyNJfOUgZTBPnMW13IEKvFf17q76iqS/1EHm999qWD1x8CaGc4FTQK2/mFPgFAfHqzRL
MCYP7Wm7c3kokJZqlmMZyMtQDEkVrzKW+89TKhuKb8YzzGXxN2Yt+imtwDQjGBSo+wWdCClWAs/V
yCFhIBbUbgedceG5OwBUGPzF3cKFdfTbj/fYgxu9nBe0TXMouJHTpodNNRc9X2T0+Zow1F8StNEA
DfUwLgQQTNDsmuTiAZw3Rc3WP+E63GHuZIioZckyy5Tte+pKPnYB5JuuAiYvHa+2BiBW7mUvaI5O
Hw1I5uTWQZ9uh3q5zf1dAaPYOsSWenXg+gHNdnHRQe4jIpZqV3sg6Y4LPysOixODsfFP2VgotmgN
PMZIJWHyacnv1YFx2e9RL3xYqJI7uxsK6XJrjzSp4X1JqwwewtWJHE12uPdicE4HT14VNBwxylxA
kafq04UFOqRb2pc+e378ooFj8gFNWLJIn6vXUSQ/v46IaCT1qf8tkIlkQwve6MnOX9JSDJtHuJoD
9nOeNWJE8rHBjS2tY5/WhTEJYAwHe2p7438qT/GK8D8jYguE7xTh7dmU+A2aPeYnllSbstXPLqo6
bzkE75gW7udORP1jREsAhutsbPeg/zUNtYiDZ75fJE6JV69UAo8D1OHDt0m8zD60O0CIVE8i4HjR
oKNUpZ/lx+V+4v8RBEb0HeFME171DRhJ5mbKWgozX3kJ96DRuAAUJ8oOFDuC1cze8dcKWzIfbyka
itDxOEjRMI2uD0L9ooMhguPjw9Vecih0hUww4VQkJDkaI1dxgG/Nq0/Wf6BAfSlFp6dF4u5dKEYY
QMUrwo5QSkoGbXa5sY8FLKRltp9IssmsBn/hL8ibYyqp30el6avlTCHlCO3/PhMYsjmWfJFh0dWp
otm/f63x+9nMxoLRwwCIpzvHKBV9gIClv9IO2yPP+LCmAwkCf3PyhwaAUM+9JrvOb3Ff0nPwaktg
3rYKxHmBAd7VBYvegfO+ItxuEmYiiwbE1cemHlal6tVJuM+wJo3h/Snjgpe/Eg7/2AaMjdcWTZeW
RuigTZ/m0GjnTwLIHboqkA8nVdzeRGnQGQJaDIzH/e6K8JTWmtWkjaqzkU8WaaQfu6+OD+VmuPtj
LFM5SNL5zydYiA7jhREWHBUvnamORAVQE+N2Li53rYbGQfowtcPqc0htOsjDQ6fFH7CxlSRz0uln
gDQWAehEdejm/5eT+9DAU9tbo96NWB6yR4el3EMvgWVTxxRYuj2Yd6CfLeW0WE9SA8EyPVExD++a
e2aEY7cXO6Gy4cSnGRHoLNAdyAwWeFOQO1k3sAtVL0G1IBhAhV8rrUP7wE2w6WeIaDtsB6IPMKHf
m4hRIv1ypqs+0bvbnOipE7/5a0AQqpmqy7n7ZBHSrvxqAK0jz4sSHEKU8DN2PvowKw332KbN4tWw
x7iaKQlTax15HAHHH30Mw2Iw+cuA8x/euhEOWudpc2lkEM7maWmdSQC93RJrNI+kr7iLNVsFjoKs
Gnl+BeyZfaG+sfQ1Hnw/T/FGdis6U8td3C4kjgfV1RsmrxaOzK+5qwFboiAxCopJW0xKIs6R8y6X
cYM7u1Oc7neTq1PDmtGhmchY2d/OSNy+i0AB833bhYwTNbxieCS8eikk+OmXhWvGmr3rIAiCKEHQ
uKSyzAttBTeFVesBZxX0WkIo/E0QHnx4lFigvzbuPRl+X+Lf1PfrnOjooTSDuv7Ec6zdmrTJHPdm
sl/vES8h6oeP53qcvqN0VdlZfyk2ApZWyDB2O3jxxdWYFAq1/Q07IYJX7amg+VBJZ3r8Q9tGM/AU
bhJ6XecCXt8T/Dfe4WSTUGQZHBGv0GFm97JcT/j10rJqezeU4YxntSARvf45aODiN3MKXE58CgWR
nwDyoJzJqKmkaYeFeMULC6Wjq6plV1hh1EjlBnkuYrWvbxox+Ku3cCxuE1TiH623tcNarINuQDfb
z8Xm97RHlc10+MI8S5iCCiuyUsVBg2qCtxWN+fpteB9Ur7c8YSTAIynNGI6LXVW+AH6148ZniJJ/
o/JcL+IJnbNpl9putKBKGiEZNLi3uV1IzTkPE9jRSXuniCJbBwSQjY5VRx/dmW1Umv06ZCdTlRvp
HuJgxho72m+9RoHIz05HvN6jAHCSLNajMTdLGk5zIthf1nni/k/q7H9u/XEqxliVX8rrCk+1NMw5
QMiauxYwpDLTbv6BBUVWDpjp5eVT0Opnd58tnjxAdPvCsKDl1UnZ5fQc3cX6o4if/8cGPOlaNhlh
cIkR/CZ7I30p1+h5Oc6Wj3AHDEdfVQL5m9EL9yCkLl51FRFSitOAUxxDM0bu0UQM3oeFDvV5Gp7r
kgqzPUCEQVTdG3hDDZ/4osAkEjV6w//4a+2AKpDR6lpfHRoistnv0tujgvYzm576dcQnnzJzRbjY
B52ZkQSLQqhmCB6FsYqsAvNbYLSkK/ycEbbwROdX7nIqfjRaW57T7WqKF7VxKm74ckzzDCTmF0hc
xPZtwSj6mgq0ng7wwdSj5gM98kwtFcCmEhVyyDbHUiuB6nBkbrsLXZjgqqRTTe86iNmvgvZz+Ayw
h/i3mm6M6lHEgzSe+yhueqBD/rs1APvx99IvQqBGZ1WtLAhfJliTIeEO8aMYExbID9tlK8wyb2gs
RYMKrVfwk/QPB2UNmd2nzh+GOaBrxi4ytmc7mxK+sAl7IxCO9+C+ucH1dVuelYx0gMrMUVL7Eq1d
oXOIT5d5o0NSNQrbI3zPnhRJ0LaRbVoPPtchPDxTqNpT+n+8hjSZXpc1gREANzjqvp/VSBmk2Z/M
xTARqZHLL7ivyqX9RfSTQS12/2wVd8MPgbtTAMiWNohRxdWTp78ScRuVzAjbMOrUd16kFTlS9Of/
Vwida2NBXXUOA9uwYAUggqWUo/k2jGJVsdamk1qoVPQswCO5FkFQMXBzF1DJJmVdHc6AAOAH1MX9
eBuuAQrwB/Mnw9RxxUaV9otnuxCvGgMn1qmnsjM/nMyNT8bj1TrzhG5P5K2hHM3xQfHA2MDJQtKf
Fp5a3n2bAHhTBRBN12TcbpBelxuC7Brm6Ts4wqG6QzG7NZAozT31sBPsrkpzR9zJZAIsfuxAr6f9
TzIva/9/T6OJnswaOE8XyhcyxsbAXD0byxm7iVTeMwyn2DoWdZ+rzVS/fqLLFSqJY3+4aWKQ9pzZ
+j0uBLDv1Sd9GxiCr0v4KKipPUo7qJ/3WikqOQ2jNvsxs/2r5ccktGu2/C1RJVDNy5RMfiCOud+A
qn9zmqhvmvdHigQIs0mOWPiR4yDmb6oCaBE1pVVvWkHG9siED5x9PCKlqiy1WlzIjmnbO6nL/IvL
ANVKGkKb3SgfDUOVDYR5VVvUJBVLgvJzbVXKlvRU5TMRza7P9gKCgWF03JyvkJ4Ko4GUoQ5abqA3
SjxSCxtqszmT9sIoNnKS5aLfRsZScsBECdDhA61dVrwy6n1HB3mtoZ3QeFV7ZX74P11McPuHyB3T
1nqEZtyQ92ThgcAFocexFF98/EnJRg7QL4ofwhUB0NSUycO34il69cOJDF9h2J1WJRmeDkukn2AR
xUVNtpW6s5WIEiKeBJDOI6tA3Oe6wdvS/8qNeQ4i+U6OOABZ5KQ7MQpeDjTp2z6bmy0xBltcMzq5
0PvZwmsxtTW6GOges0USUcovTHPxazvPHsaLKEoyO+uUyTKPoRxCIcut9FuopmhgX2b2yl6X6SGS
+4Vnof7UM1F6QHOWiTgx+TfdEcjE6f9im6UhnzNxCswv7nPOUIdMR5PPTnJeYc3AlkE2Yjk49BV5
7hrBYvBGAnImZ2PblNSR/vqJDuTw+RzxLY9vX709hNhBiPdehmg+eQhxysxJNYy6SvqdtTtZVdzk
3W39bv5ctKjLAJeiDGbg8M8BSKJCtY3kwqeF5rBC2giatZ9JeuwrCfolE8vVFQiwCTQS3XjNbalr
Yy57ULVhTSe81txzecix+5n6XX3/qYTMAVfGfrC3mnszG3QThJCuxDDYv41LNHx2eNOceGAeRpWl
A4vuADuHGFS93breBvPDejDgdryhvX5WgmG6Qdv1jz09HVuRXA3iQafj6qZbg1haUPfHmecT1kPj
Z0thE8gNzV4XcR+IXtPYGzRqDk2/29j+t1JFYPBAsG8LNl4XoxrBw1gfUGJGqUz9zAhrKN7ZDZpZ
DmgodxVdXzgolCTV12JqHBdGhHiR8ByLh53WPo+DxnJD5DxB35rTTXSrjX7oBreMoPR3yqjpx8am
QNdPEyq8E9aOAqtNs/LXr3okd7zw57O/Vz27nKoAbBE9xndmL2t63Ce0WBhqtrap5tZLZ/89yT+X
ABT1EJtxRktERo4tZJafbdMYOv64VXsMYCCkzz/zn0/OlE78drcxfvBLs5aW9zN56MxUJr8YZX1t
F4dK27a7psQHD+HFG8+MqHFSvFA+bqLK+Nr05XyTCWz4TQlfxlkFOLJKXqVG1WUybTs7k4gOuAVr
b8wRVonGdK+6l5oTAKV4CJqe3f6TeRarMTBmn1+DWlDmX4CiJEQqthIXFyyVhIsnU9EdLJvhrT3A
J1SY5kk1qTNeOhXPbm0GD3AAytDDHBwNQRth+YIlMW+H6pLVyO9w69aKYaVcprOUFE711Bg/+jVP
smQfROGgghSN2ISsuy4T9YvPT7q/UysqGiBIAxtzmMkK8jadx0JiaeW0rNdMBdUrI+WNaDcD+5UG
rvfEmRbfwmOAPW5qp6Dc8zr/Zbr5oRh/cvC4xc0KI0eCUmyZp//j5foWwhbDW08SMYzv2bDSR26j
f9LLiP8m6ZDxu6iCRbYTwdHMhJa7oWQX1vgWzc36wTD1AGqu+gxQUzw2zfXNLIuhEyvgU8q3X0O+
8HK7Z+ghFnwWMppfKimO74mydq0USozcp8QyIocJ9kVzqCAG4M3sTZEFSaZ3VeR66ajuQDZhd/b1
1/tAMnMLUBHlBBgMn1qqEpDwysIIuQSqgrxOmzZBRFg9uQ6g65xiKvS6/T3ey9rRww0Bl+My2WKd
4frNMstIp1T6ynlkI1sw0q9IIiKd5GfNFd7FXF4SGiMABeWN2V+QdmxehW0x9WjsuDDzsxN2Xu85
zKXULkhcKJ1sF9JNld1f3PeDzdw/PjnlgMywV/KC3IBdvqiQlkBe9nECfuTMprKVT+UuwaWMikl9
JYHfhxZ6iWP+Cged2fp1IRg8cXEgeVSY9RhBW0aSgsXmlvEddbeqSqMNqRPIXJkjYdphE5nEIoWq
FA6YAVkCkCbsy7/9izHcVXaIY8vuNoad2aaCSt4PpIkhtarLGUBw63Yl/9vwZEoMdPyvzvgIhSLR
q0unY0yQ0V/J90iPx03SkeMdrrYUCr7Ou2LL++vaym/Qs2QCPHP3YgecOWLCBPMaXcLscR/d07yA
4GKVXf+RcZvrbZPI2MR/P4XfTZMb9d/8/N8qoIg3EDlk28yl8UnG4EhTd3HtUQXPwihZcGNmnAP4
dIxj0BwJoRb4YpVD8QEILwOLNSkbKmXUtfOz9xkfnM9kemcqbcIB6MNqsTfUyX+HYzDFMY9XUup5
zIcrk1ae4wZgf0pb2OYYWz+8wuTCN4l5OIWHG4p+dCehm2qvpX6SvDmpBGXyTT2r6DpQVVBcaJuH
Tv0IGZ+mZNOxi8mKjhjR7Iqvs46Mg6zTdtCzmCxXDjGBr/rZqYMZW3LrC/c/QuuCbsE7+k1/ZTd0
CBD1ulxnw2kWkL+NRxdAcIXEll8cc2G//nNW6xIYEaToxBop9VhJP+SQ18uaZOYrzsD8WvtSYMp6
HVIoWgEFGvQ9X8ViUWquIh4pMbfhFU5UP/gEaM/EUjeytoOdcqhmg1fehkYBh0x4LrOvUUI+byuY
g2pA4sY4Tsg15qB1WCOzK/YZHR1lRX37UA14pdSq9ynFDzeGQ/JjDCzbL/dye9UJxB1Rh1ImwwEE
G6+3ZmacWs82IW5u/iBpzngCAfiwxMKlXaiGVYOAlewy6+cSuPwgGrDFXN3FSkxUWCgATUtRLEQE
MpTCl+s1QIRCd2AE99VIuy3SEahRX6+hyb0U4Fl+q/skFr4Cgm9AhagD8i+qnWlkjqfYS5iEQYBV
dn96MeuFtMUEx5zq8UCse4aBjOh/q5Q1+Z9vQUgzu5rVW9KJpzteja9Dy8EvPaXZBx4GjkznD1CV
Tcfmn6Wd6PwsvI4lUQIb32k0f0vUozZpvOP2yfy9buHE3ZUmNfXMow6vpjALpeAUF+xhvJuuacXb
5WvEvoQovRGd1otQidI1pd9FqB1s5IceMIIDzhdmx9tkRAaGsujA0RTFzsBmUGPTwVr4EYZ+ye+O
UbifTLBK78OSYhsmzPJE/UVNCQsW5CBbQEGdS8crLix0gi6gyrRtSu+tUDbY3B2DcYqrEvfr2xwG
pRQCx44ZKaA8y8aKMfuq3Ffmt3g8MMkIjHaz1WYLlwwDHAmQ8MymFzVQemaplBZSnGNdTuMOfo3O
sLSvWse2sRVnqcPJmtZ5Foyb3InjYeHzgdIdC/n/lFVaeceomqyx+82v6+k+uKjWm8jmmxat/IAz
4iXJ8tyIC60VuCsCvgDjb8jsYMD21cVWH6M2OKbgt1itU8Cnwz5zNqR93CmizK5MVkGbhQeWpym0
JEEjkW/pBRi/LhiY9iJB2qXmlmPAfNurBbDjdC21eKqzHtIaOp8duHl/mm+l8RKGb6gyl2QDHLD7
5yBDh2/0HAj9nlTqejgOqDrJVWdisWfkQUBHfds35KS9QeNwIcw4B9V/S8Es7rkQyI49hByqsxUl
3ahlfKM2S+07feoRxJFPNHtm0G+v0Ms7XtVfZFrSX2tFlQDCtAvmCkHwicQwTdL4KBXCjwRKpK8a
8BD5RkTuYnpg7VevXLXUlXaQmItYHU460ORh6u4pdxG0P+wx5yGWKFpXLJS3DjxcJzJv2S/6rhEA
2ca61hCNOXEjMc+sVgvgoiWanXu7zjVeXKN+4UsxhkK9qNLBST6Y5ybPtnweksJLB0hx8ofxZghu
sEW3ZWIvuOOteNpY4j9NfOYQ22B9WgDBzn5bEUuNC4U5TslZpV+BR5G9stlVMCuMxHE2qd5FJ9bM
Vd+PVXCg9LDJJsAD3oHNAwoHtdxKRijRyp8HFUe59jK8V2akNz3xD5rruGHEjHAiTIwEDUKBuiE6
CkJKTWxyOOkvN+/0GQ+7G0c6lxAbF1MC9rSZzARJi1lp2tWRQjkKA4Pmfi3FC6QUiPQEsR7DSrh3
CfjvCAbDkV7vvSnCQeQ4ahxhIgscf597JyxZ5Tptmsi5Ebftj5SVomotMLf9iDoViebRHxBJ0gB6
rpPTN2bFMbQ/WVbTC0hF1ea7wLSK7cRuHR++TsG4H9LRVe/IK4nqT50Au2ypj/F59ooxPLXO0Zb8
0ZLpFa7lWggCjpha8e6YA6MZuVmUck8NShCQqJ/1ve5Ab8lGVozvJs12HXaoGow3tvYZBC6I4eT5
+/C1465KsqxOcJhzWss8nICZScMwVDJFkqztwL/pF3itwt4ppV2DOumHcdtXkMBh+jCQWfOy2gJd
yYZfD0lh9iGVUF4+Vojeb1hnKFcxlCb6qApGiEf9e1KOZkokqzodi8Al9vfL2NRz9WueiPQzEE8X
VRZmbN4An0yPBx2dvL9DecYTo6t/H9I0g+w9gSD3unvHhX7khpx+TSNnQMgUJTX46zjCeL00rWYI
UlnSk9WI/dzzk0Yys6qBzxWKp8wWe/l47ffzELdgM9RffnsoG/i/zCQK+YlpxIgIJds+rB8jowHq
6P0WwptgBMKLgiTxtGbn2kb4r8R4A74qjb4d+mJNY40zN6TLS3px1gp3FtM2sdmSxLwlHC6lhhMw
SNmwaLEvRefGvRL9vHYZ64nMCBC29djgVCbktnht7gc0KKjzV6OwJqeSucy5YWGW3Fk2RDm3K0DC
DOrdRRDmfdL/m3mwcRBRuPu3sPGHM2loLR+szJamHaxxs59A4qBG8m3leVS9wmpB+PKv3RN4Whev
OpQDzU03AdVbobR+jCpvz51jIwT+YT8EMSKNABs2fNmucA/0RvqlTuFG56wxyAP5MWqMPflY/3TA
96c3PWj19NJL3eZJalOAuqCBQlLapdlxmPkKmRItK2wfTUG0RMP6WT0ld/faMFvGeaRj7j06N+Z0
ewRZ2uZXACHcm8jd7/JO+Rj0xTVUo3uLOlYLRIu/rfnJUf6Z9xTJbYLyqGDHmTzTPmAyrk5XAhlI
aQusmRv4wQnm+2sJ7lIWZQPtDCoa6XiIx2l9KnXMJSeHHYlR9YCJmpg/FLc3bNzezBYVA9pjMkpj
g+6qDae0KIbVcnc8A2UaTtc4FFxIdGUjwcsP5hpBrP72PObHsOHdtqy2bGjR9NQWtkAcVrTwyc6C
kfVsscLqJSjj8/NdQGVczR22AaXnmy7TDqwHWnUhUr6hjbI5a0878Ne0Fdvy2cWXoKhZr3BSryy0
A6PfAbAPfcOlh6sGqjAl2g0k33Bk48wlAWN7LL1mn5KYmT6QxtQKUNAk3VIaK/1r8tP5uwSoQnDF
CiFVWxEpxz1mIW1dJvxBomwMzVOUMwapCmY+RMB0NhnxXouoMLxCNQO2vbD96lA7YQ8+ybiO2nPt
S8YGrcgRytc2q3CTv2LKdlnjavX+Vph8e9csRQ9kd3vpL9Iouj/x9kh/IEAqRZVdZdEN/clhZ2F+
S7dJhgEwbI16h6k5NQpqnJrCsO3YZPRTBXFdKvUoj/YtZx6mJWW4VsYnCZPAqBtwGT+5AYUQevnN
jz0xxdwP37iabp1Qw++JWCrsmRCKjbkMLHa+i80dBy168CJJnu5/1I1n2D9wPeVnsXTKhnxG/1qf
RCG7mGurMJDbzqCgKa9opg58GrvPS1Cgdyrvg8kcNdthC9sEsx6sipMMGO6UaBpNEMyvCEVer0jp
H/kgd4aSNyUyx9nFaF58Y9z+bksXqH23l1thIlsWeEdutAFrv0ZX+Cp/CU+Xh4EYo3oQ4a6tnftX
3iCQH8kH9ioPTABNDdnMG5OSkLE293Q9uQAIvHOGSZ4awkRJz+UijhmCWgDBSqqCNKwg5uNsMJT+
2b8UgKaVfEUfrt+aQa3TVSvucU/+XREBtJvbbm68QEOYIcN0AZw5tFwKDIWPOcEhDlg6VQtres4z
gx4+GNSGhR67EM2qcyMnnGfs0p7FplOxySf/rcut+/VP4yMZxr73NcjW0pC2ia0f8587nE1F+Izm
ZRSrvTHkVa3N14rRQQkG75dTRldx7Jnf44RguzncbZjY1W+IHbD65+F+1vDMolJxZ7RQozj9h48Q
ysOiHlXdw/QiSbFG2duWoMCW/rdwS59nRxSksjarTRwtezzdaynmvfVuRo0Z4D8WKzH4ymvmUsLF
VE1VUV+5WndfHHuV5okwSkCT+2I1mP4tXTT5eFHFPmyq+Y6AZg9Six09mhOyUxJIVhtOdun47aHP
6WoLsVPpIoI1gH/WaT0HPfnmbckmgvNXnlZxrdJFa7TDKDgCx+7u/6nnbitgA3ZZu6MnDXXIg3P4
zWHDs42myTbSkBAn4/kALEpQibUMQz5nPZFFiAwhDnlK4NDF2CrCSv5Qn2JcuxIvzagj9lP0JDce
eirdW5urmX2ijGeDfpoKVF6obTwX26mhSpGIe2FbmRBAb2Xuh6zQnNSte6keowdUXQXYlLpQ4KoV
u6HxWpO66Vabo24OndA8Z4aFeZAE3kjLKzSLJ5X6UQLeoRVG1qYDUdgDCB54lSq3bGApdaYciuBX
YJ1ZLDxTL6yaVmbOeuRdOF5j/JrC1LmjxRMhJxr14hM11ojFoE3i6FHHcCeuKf4DStOnTa3qRlZ7
AKQ0OCTMj3txr2eYsTbJWNcPIoKxi5VchzSK0dY6gxoS3o2qztuzvhdDJD+qWZOYySQ+0CnB8a8E
Pb8hVDHCCGoS17AryIqgdBayDDwCXquzugo5FgzZUjgfBKx6Gs5pHLvwDwm5WtETC8+SpdX34BnU
5c5pMaZxvMjvZk7vhuO0qnGRM2PpBmrTm7m33yCJCx1fP8S3NJFx9RuagIB3+9I7LtIjfFob97CQ
gAfoEWqaAWZH1l2d6QKpkOMcSJs7mZLkiatcWoJ5HeRuOKZxkq9ps0Lp6j+ebITXO+YtXcw99cOU
bOHm39cAVcEOFjiZ8Y3qaT5nnzLUAQ4gVUVMJe7uksSQDt7y1hmTTvrqJMVv3xesoB7JEpdg4GmH
MKwokgKZqa8nnqaiLtvkAndLkdKGWMEimSILUQYcCOa5rHB4J/5Xv2aHdc5psptNvQ2t/7Hw2Q42
PDxbZnHysLwTH9tsXDqAm3ysUBRJ+AuaQ82plM8bj4bpF1ZiLSBugslfrA2KFYZNwuUHEYeDbcPu
XtZ5jneOVHRbfbD7DoeGGlhXbaZnKeq3QORb97v9T/m9WRwVkUxDdecI3yvwy1mybQeasdJxMIpj
fGLZ6p6aK5f7ZztmwnSH2mDdH9i8qD5OWd9/bvrDPodVhypApAXW51/dgYln0qO/GEEPM6JHeRZN
WQ5rqnu+PzRHdpfiPcaFqurP0GmiJ6ZmuN8zwldZ//gycJQQsW8B3zP7+BvWALBYXsr6fUvUoEUP
Y1lbvaVYTbyRj+GSbk+MoaboeV5qFZo5isJbe22wc6tbg5+5C08hOoAFuBnlO148eBuTrbZReI2/
L01+gsLaP0IAMzsHvUTt0TlPhvzSKrdE8tn4JezHuwunvCfYRQuOwG/yoWTtvfu+mGlvg4kn+7gF
PoTNwUdHYi2jkoCQtfjD1uwsQqlPldYE7rYNE9/nZn+fWm/sxfZsxj0mdkMeKIdzPVT3Nfe/rO+7
lBeCHvWLr5Y1yf1GU5hiZdVCsJNLH/IOVS1iEo3dF6mOjx+S8EafXJ9MEHCDp/+S5nFw8vgivZvG
+3XMGyULTyvQkbTUjTQWBmfeqr2H/HJt37KhbO2s+dm4dQCygUNkR/UZlMWl0uJVz1zNPQsuK7I/
N4Rzal22SdCKcx68rJ73kYZpWR6T8i5bQdAhmzydl0uRSASnhp56vQrzABvpnqjqEtrqB3DIE1XM
R4TzUgbQCSogO+pVwpGZIRoqKhFvcTpYTYjfAGjHw85boz35zaanbmROsmfxplWScr3shtqv88oC
NP2N1RTRonEc2+sfWYVGQO69e0BSFtFZC++tel9mFZY+BxuY8Tgs/vwY3tRgXZOOxaozg0s5bKKn
2U4G/5IpAbweaoefBR3Le20YVoxofoXuWCSFkw9E75H/XEHoEyyqQ/Mn5eIdBX9Iw1yFYMW0wYba
enARh8192csVYDJaK3hOJUUaw+RWhrwCwImryxBgosm21JOVu4QhTaqWU6bayMZbpZPnldt7ozJt
YAcH2XE4H1ZAjVs5KQV99jDgHC+WCNSxt+K/7ignyDyWgGZd/+bJqFQtPS0HlK/e/XS1WdJHPdYB
Pckz/ngIYpEHAkPuGubx33IGDlSDMbFEmwNnG9c4OKd01AM5KfyvzzqZIv8Y3QFwbvxWMpc6KIB/
vUQ6XQ8ISp8sDOEJ2k62Y45FAY8Vg55bLzaKr3G2DuWXDeZO8ZRwHl+IljEyTBb64j1Z0Of+Nmbi
UfIj4OjQ391YCLlMBk1FOdJ15zxZY4MGx/yd7qAlF8mJHkMZI65zKtd9SwoGsVpjEauIS/6Bim0y
MMV8/Cl/9jQlMdZI9ChXX3j5v4e+xCvyRcfbG+vDwU0IlTQrU4+ZBq0+TvfKz0ocQT8AngxDBOMv
qUjgOlBt3lWaYfbmlT0htNMw2bvuY2tgzsgeS72tevjPV21WDh42j/RHli2Bd/5OEzstBsvj9Jxw
FFfgHPI24oZ6M+i//vOJTZ18leorknQwPhReUX7tR8I97pW2+6n7JG300ivtVi5eQBoWYyFWbS0s
vKNLIGm2lLjhdNDrr6+ZsMdT0ttm60iBO0Gkxr2Cpw0oDY9TExK9r2HpTkmgPbxODH0YPenc5Mhp
kE6NaPzMWBO5DPL5I2hbUS+foHWc0km162RZoQYZsd+20SwNTAW5y/4ChpWjZJB7Japbd1t3JmZi
NCFIIAlSdCo2h8UIZSQ0qvpvcxfrUL1o+blJv82TIMwA7g//4VPz7ADH+7F6HOFW+YB2uGQGEcp6
t5z3gI7pMxx42JicfwSDA2bEw/aSQtKvMcFWIBqHTw6VRVDvr74l04F7qSSYtrUi5lwsosU+b5BV
eNReUa+nZIQMX7j0CmjWspWgoxmb2P/goiAzcJDex51XL0Uv3Qfp2squAEPPznhoYnJYPKTn86/9
BLndFz7OR2usBGkmKFjKHEorQekHrr1bOUUFWcsVyiu/G/ftoCjUZvDmeSKB0OFvBzKNRYYpDKpY
VlEw0+p8Uye+fsGw/VwlLYAI2Md0EH6ZltlfLXlM9ctwxJzsG2YbPF99gDi9lYxtCv9Y/oX/P9kH
QK3/yHYCdMA2isFiS76/8wsKBoLBexV5VEzK3+tYZlW6FlS4LIdh/g85sYohK267ryTkVmwOAPko
O0uGnXqNRfDNib1ylhBNxf2dDd6Yt7OxgbojIttd25AY6wObEJNxwDwD+DOzDPJTEV6/FbpDa30F
cjsRpx4hs7/Ej7iP5X28PO/0AZP9ERXee6dfG+XQCKIZKcK+KQ5DB3X4gw6wXbEpQXB1Kg2mFLNJ
NCBFEViXeob/x2EPp92o/ESg7ZH0IEhE2ESz7fIqcMBrR0ZxGR+YkCHq5XRc8zWKGeQiIIV8BCY0
8YFimfNLFbu6IkHMvWcxmjXWEfB4enX1s5wLz8lHUSEzv4v3/JfRT90DclGujrQnz7GhZ1c9khsH
yK8OQwlI1By4BnHuj78JQiX1hXqLdAbkCMLhmf+V3g2eLxVBJ4mgsivbtl5NcOVMJ7C1k3aGKgHz
7SZawVCdupHSzXgAxmRUwTYwBA8irk8Oh65I19B4mIzRP//4zYyGF2iDIyckbNU7a3f7ccC4h8j8
DxXxH9lQNmOIPWNVAN8TTMHbsUb8AaHixLrxj0D6B73XwqKeKqPisXjd17Ik91Pc/2tEiYcU6DtG
pfKKP1EAHGEaz+YXeVMLyGpJXYeiHe60CCH6lQIczlU2ag0692B499ENoqGbfoiZoa1iwnxF3ugk
gmQFO0QXvNZ5r7FVPZDk7pnQKd1Z3yBIjG3Eob6ofDDKmHeAlkAXjiprRD6QXLdl+F8ntLzDfa/E
2IeNwJdsrjQUOZZauGIohdfY6hbQfqHTWgwJlCcmB6s3xMkl7VwYLNftBIgh7DJ7jC6CLlnI6kpp
ojzTmtMm4dgwU6f/ZKnqYaAByzjyXCkiefbQVKRP/JkChHkOOAsANzC+fydmqoHTz2QmUXdmDL5O
GNc6/NJthGBqzpeCco8gbwI587vTxFW2uz3RklgBhRCK5M4xiull+4hz2fQdQhhVIY3ShChWJMWc
udR9LrlH83PO97LKus+bIyDNlajONvmF+tN6ibkFWcpwwSBqjqsnjyDwxYukfmNfPd0uQ+eREp2F
Gg8uHrfR7Iw37DiCtv5Pa1OjmY6Ei0tSlAdSvQ0S74TAIY1K4DTkZBWv5nxzur38Bhnn436xANrG
M/5W12DyJCHIjnbaH//ltqOSayH2mBX1ZTFZCoRaG3ZGdw/1gkpC7XcE6D40CEKxztnPxsA7+Y5b
jyXBL3Z8OK2Bu9YklS6GmXmbICVRP11prupQWSHhKhRhbroqEFXeIJcJXgGevuP24U1qAt+oTbsU
2B1b7D5SibXMQNgMoKN4t8Q2Za1wkcB8r8hGmmu1U2QG8nUyePvcI5DjcIX1qaQfp82C+4IoPYwy
YjXlVckN96rBIookImL4vmZgOMve29Ce/FOLgM0yfW34lICNIpxrafg+PSHkAYMrWP+TojCpd48I
/8yQQefYIf5jv5Txw/s2g+70E+LPIJo6ObbwIslOhkQgbVzOBasUspMcOacOZdgxWMFte0/9EAkE
//Oqx6d3Phd76/aD1X3yERMG//L/C0U0qsbSuRbe9rXlA68dVPhlnYWkeKOgeqkYvqUNxa/nTVKz
zbd0tckr2eq9/2mf8Zt9w6ReE+hNkx3RsGCpWFh/RxO2ysvVyFKXRC9nW0Z3lVsqW3rCkPVfbNd3
rLt7o2Lx4tPqHqQLdezTV0CteDPMRyuzZYgGQtCww2Xu26uThxMjxLkd50CbjP45elgg42vHgYBh
4oGhjKoZksrPt7VYbaKok9t2PZ5AxpcTRTzL4ldazMjALuhOlpXbLfVuVF19sy111H4PfIZfCsDk
SJc/WOH8fcMcV8cehUsF8aGjLH0suCmCkzC7MoMyCjPoRZKJHhBbj/wfdHVwiWK5QL6YSNsz6rgH
JBOnKg89XXGmOXdz5bmOuAAhh9yFZO+dDxbM+Kx3ghcAwuU2eOXE2piZpspCj4TXMUSfVNeJwo8l
kCRSFALUfCipUxWSNYg3hWPvfGvSxRvTA877JBfcQAx84vf+AofPryvd26VeScF+cKPNDz3BxMVK
235O1oS4VgTShOAhQ/6ku5DaQD6l0ZMEYH2MjJkXc7VFLf0qRIQcYw+vBZ5WFvIJ//QapMzAoznO
nig2dreKGPlf42+8nNcMPCeMQehu2EQtPaH86An1Yk0yobMpznljZfxACRu8fYQ2QBllG/QqV6k7
jAKpOScxjuuDSm9Zt+4HPbz6A5/z63XeZgoB9+9OBX8pe9cA7wCcRvr52drFs8geUIWz944K1BXC
JlBxSsFMrN9D8qQLZLA8iYdRkzDYFbMh8yCXuFjBXt2W4kZVexT5SSDReEVVHH/CrgCAP+zd6O+N
9yj5WMK7j78gb0a8MmKBPL0W7gQI7S0EXkvJP15JXibTB28hcWsJCj22dOvREd2vg8mj660FzAxH
u95uU21WN38TSU1O7+tsCUlI+Tv3Y4Wger1yzrjXVCDpzUpbYFuALXoNZO7bxFkqQP9vPYvPbVlm
khmKxh4ViCYUyFr54PfWsEpPtZx7jgpJb1lMHbO9gNf4bwImmP40fGlmJ+DI/7Yb0dLJavRp5Qyk
SIQDwE9drvMvuDMuZAgBGGjhFHEthuyvzKqGGJQ/I+bmg0rCGZmpwbvUhVNdNgxd96OfL0I9UNrt
Qu4AlSpel2+/6deVNSImemkOYLdqqrfj1B5F8fIu4Zjh8suhP449JXYM+9sCwUiEcitf7gldqoGr
wQPsDzsgTIOt/uhYGr9AWa4zawXdDipT9pg6pFsxXJC1nQVbFUc8kKX7dPTQVfek8HdM5FAtWCgm
TaEHZQA9BArUDTg6sUlQTSOyYY6LwZWgb1nHgoK56xh6ZZQMBFJw7pn8w1J6C75fcoSD4ev7TIZo
/8BkU2Ah31QKWIfUDhr8TWaqKLazCFD3KfFk/4YwozgZg3Q9UGgbCpp0uBwaOdKDq0RijY/tFUBa
uYpKWkWcv3VzfY19B/YBJZhTCaRaJP+NBVKJv7AazObXK2xApyqL9E7YmoP+V9XJ4p4r8lPbG6bp
iCpNaDGHCXXcUdAr/ORGHa+DpxbaEO8BM4LtKbqA/rdw4ajnhWYoUMNn0gFtZ1vbLsWygfLSQoqe
SXpU7tP0OzKAX/ITAN5bob9NopBb6oJuNXdUXtCXbOSQC4+Fcu1pUIo/9wRUhVDBg1eKARWBmX1r
6Re3W1zl/wMFbK3A7srT7Bqbq6AuBrlVYIriDASMNppjOEjtF9q7yaBkmhODpDYVlPtO1qcbwQE8
5d+JkdgynZatip6E7rVbOAomVZI2398fuVtmI+Qh/8+Tf/V9PC1GvMuXrbVPWWARvK9FTD6UL4pE
/L17T5TN7snh4vzxQHK4h8Kzb/2OrUcuI2Y2Ymd0iQOidW/7RAQEMSeul5l5gDz0Q+s2RUu9/zbx
S8msbes3D4VLr0AMktS5lpLsrJvgL8nmn4eVHmsUsb83
`pragma protect end_protected
