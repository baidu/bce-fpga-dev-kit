        `ifdef USE_DDR4_C0
        .C0_DDR4_act_n(C0_DDR4_act_n),
        .C0_DDR4_adr(C0_DDR4_adr),
        .C0_DDR4_ba(C0_DDR4_ba),
        .C0_DDR4_bg(C0_DDR4_bg),
        .C0_DDR4_ck_c(C0_DDR4_ck_c),
        .C0_DDR4_ck_t(C0_DDR4_ck_t),
        .C0_DDR4_cke(C0_DDR4_cke),
        .C0_DDR4_cs_n(C0_DDR4_cs_n),
        .C0_DDR4_dm_n(C0_DDR4_dm_n),
        .C0_DDR4_dq(C0_DDR4_dq),
        .C0_DDR4_dqs_c(C0_DDR4_dqs_c),
        .C0_DDR4_dqs_t(C0_DDR4_dqs_t),
        .C0_DDR4_odt(C0_DDR4_odt),
        .C0_DDR4_reset_n(C0_DDR4_reset_n),
        .C0_SYS_CLK_clk_n(C0_SYS_CLK_clk_n),
        .C0_SYS_CLK_clk_p(C0_SYS_CLK_clk_p),
        `endif

        `ifdef USE_DDR4_C1
        .C1_DDR4_act_n(C1_DDR4_act_n),
        .C1_DDR4_adr(C1_DDR4_adr),
        .C1_DDR4_ba(C1_DDR4_ba),
        .C1_DDR4_bg(C1_DDR4_bg),
        .C1_DDR4_ck_c(C1_DDR4_ck_c),
        .C1_DDR4_ck_t(C1_DDR4_ck_t),
        .C1_DDR4_cke(C1_DDR4_cke),
        .C1_DDR4_cs_n(C1_DDR4_cs_n),
        .C1_DDR4_dm_n(C1_DDR4_dm_n),
        .C1_DDR4_dq(C1_DDR4_dq),
        .C1_DDR4_dqs_c(C1_DDR4_dqs_c),
        .C1_DDR4_dqs_t(C1_DDR4_dqs_t),
        .C1_DDR4_odt(C1_DDR4_odt),
        .C1_DDR4_reset_n(C1_DDR4_reset_n),
        .C1_SYS_CLK_clk_n(C1_SYS_CLK_clk_n),
        .C1_SYS_CLK_clk_p(C1_SYS_CLK_clk_p),
        `endif

        `ifdef USE_DDR4_C2
        .C2_DDR4_act_n(C2_DDR4_act_n),
        .C2_DDR4_adr(C2_DDR4_adr),
        .C2_DDR4_ba(C2_DDR4_ba),
        .C2_DDR4_bg(C2_DDR4_bg),
        .C2_DDR4_ck_c(C2_DDR4_ck_c),
        .C2_DDR4_ck_t(C2_DDR4_ck_t),
        .C2_DDR4_cke(C2_DDR4_cke),
        .C2_DDR4_cs_n(C2_DDR4_cs_n),
        .C2_DDR4_dm_n(C2_DDR4_dm_n),
        .C2_DDR4_dq(C2_DDR4_dq),
        .C2_DDR4_dqs_c(C2_DDR4_dqs_c),
        .C2_DDR4_dqs_t(C2_DDR4_dqs_t),
        .C2_DDR4_odt(C2_DDR4_odt),
        .C2_DDR4_reset_n(C2_DDR4_reset_n),
        .C2_SYS_CLK_clk_n(C2_SYS_CLK_clk_n),
        .C2_SYS_CLK_clk_p(C2_SYS_CLK_clk_p),
        `endif

        `ifdef USE_DDR4_C3
        .C3_DDR4_act_n(C3_DDR4_act_n),
        .C3_DDR4_adr(C3_DDR4_adr),
        .C3_DDR4_ba(C3_DDR4_ba),
        .C3_DDR4_bg(C3_DDR4_bg),
        .C3_DDR4_ck_c(C3_DDR4_ck_c),
        .C3_DDR4_ck_t(C3_DDR4_ck_t),
        .C3_DDR4_cke(C3_DDR4_cke),
        .C3_DDR4_cs_n(C3_DDR4_cs_n),
        .C3_DDR4_dm_n(C3_DDR4_dm_n),
        .C3_DDR4_dq(C3_DDR4_dq),
        .C3_DDR4_dqs_c(C3_DDR4_dqs_c),
        .C3_DDR4_dqs_t(C3_DDR4_dqs_t),
        .C3_DDR4_odt(C3_DDR4_odt),
        .C3_DDR4_reset_n(C3_DDR4_reset_n),
        .C3_SYS_CLK_clk_n(C3_SYS_CLK_clk_n),
        .C3_SYS_CLK_clk_p(C3_SYS_CLK_clk_p),
        `endif
