   `ifdef USE_DDR4_C0
   .c0_ddr4_app_correct_en_i(c0_ddr4_app_correct_en_i),
   .c0_ddr4_ecc_err_addr(c0_ddr4_ecc_err_addr),
   .c0_ddr4_ecc_single(c0_ddr4_ecc_single),
   .c0_ddr4_ecc_multiple(c0_ddr4_ecc_multiple),

   .c0_ddr4_app_addr(c0_ddr4_app_addr),
   .c0_ddr4_app_cmd(c0_ddr4_app_cmd),
   .c0_ddr4_app_en(c0_ddr4_app_en),
   .c0_ddr4_app_hi_pri(c0_ddr4_app_hi_pri),
   .c0_ddr4_app_wdf_data(c0_ddr4_app_wdf_data),
   .c0_ddr4_app_wdf_end(c0_ddr4_app_wdf_end),
   .c0_ddr4_app_wdf_mask(c0_ddr4_app_wdf_mask),
   .c0_ddr4_app_wdf_wren(c0_ddr4_app_wdf_wren),
   .c0_ddr4_app_rd_data(c0_ddr4_app_rd_data),
   .c0_ddr4_app_rd_data_end(c0_ddr4_app_rd_data_end),
   .c0_ddr4_app_rd_data_valid(c0_ddr4_app_rd_data_valid),
   .c0_ddr4_app_rdy(c0_ddr4_app_rdy),
   .c0_ddr4_app_wdf_rdy(c0_ddr4_app_wdf_rdy),
   .c0_dbg_clk(c0_dbg_clk),
   .c0_dbg_bus(c0_dbg_bus),
   .c0_ddr4_ui_clk(c0_ddr4_ui_clk),
   .c0_ddr4_ui_clk_sync_rst(c0_ddr4_ui_clk_sync_rst),
   .c0_init_calib_complete(c0_init_calib_complete),
   `endif

   `ifdef USE_DDR4_C1
   .c1_ddr4_app_correct_en_i(c1_ddr4_app_correct_en_i),
   .c1_ddr4_ecc_err_addr(c1_ddr4_ecc_err_addr),
   .c1_ddr4_ecc_single(c1_ddr4_ecc_single),
   .c1_ddr4_ecc_multiple(c1_ddr4_ecc_multiple),

   .c1_ddr4_app_addr(c1_ddr4_app_addr),
   .c1_ddr4_app_cmd(c1_ddr4_app_cmd),
   .c1_ddr4_app_en(c1_ddr4_app_en),
   .c1_ddr4_app_hi_pri(c1_ddr4_app_hi_pri),
   .c1_ddr4_app_wdf_data(c1_ddr4_app_wdf_data),
   .c1_ddr4_app_wdf_end(c1_ddr4_app_wdf_end),
   .c1_ddr4_app_wdf_mask(c1_ddr4_app_wdf_mask),
   .c1_ddr4_app_wdf_wren(c1_ddr4_app_wdf_wren),
   .c1_ddr4_app_rd_data(c1_ddr4_app_rd_data),
   .c1_ddr4_app_rd_data_end(c1_ddr4_app_rd_data_end),
   .c1_ddr4_app_rd_data_valid(c1_ddr4_app_rd_data_valid),
   .c1_ddr4_app_rdy(c1_ddr4_app_rdy),
   .c1_ddr4_app_wdf_rdy(c1_ddr4_app_wdf_rdy),
   .c1_dbg_clk(c1_dbg_clk),
   .c1_dbg_bus(c1_dbg_bus),
   .c1_ddr4_ui_clk(c1_ddr4_ui_clk),
   .c1_ddr4_ui_clk_sync_rst(c1_ddr4_ui_clk_sync_rst),
   .c1_init_calib_complete(c1_init_calib_complete),
   `endif

   `ifdef USE_DDR4_C2
   .c2_ddr4_app_correct_en_i(c2_ddr4_app_correct_en_i),
   .c2_ddr4_ecc_err_addr(c2_ddr4_ecc_err_addr),
   .c2_ddr4_ecc_single(c2_ddr4_ecc_single),
   .c2_ddr4_ecc_multiple(c2_ddr4_ecc_multiple),

   .c2_ddr4_app_addr(c2_ddr4_app_addr),
   .c2_ddr4_app_cmd(c2_ddr4_app_cmd),
   .c2_ddr4_app_en(c2_ddr4_app_en),
   .c2_ddr4_app_hi_pri(c2_ddr4_app_hi_pri),
   .c2_ddr4_app_wdf_data(c2_ddr4_app_wdf_data),
   .c2_ddr4_app_wdf_end(c2_ddr4_app_wdf_end),
   .c2_ddr4_app_wdf_mask(c2_ddr4_app_wdf_mask),
   .c2_ddr4_app_wdf_wren(c2_ddr4_app_wdf_wren),
   .c2_ddr4_app_rd_data(c2_ddr4_app_rd_data),
   .c2_ddr4_app_rd_data_end(c2_ddr4_app_rd_data_end),
   .c2_ddr4_app_rd_data_valid(c2_ddr4_app_rd_data_valid),
   .c2_ddr4_app_rdy(c2_ddr4_app_rdy),
   .c2_ddr4_app_wdf_rdy(c2_ddr4_app_wdf_rdy),
   .c2_dbg_clk(c2_dbg_clk),
   .c2_dbg_bus(c2_dbg_bus),
   .c2_ddr4_ui_clk(c2_ddr4_ui_clk),
   .c2_ddr4_ui_clk_sync_rst(c2_ddr4_ui_clk_sync_rst),
   .c2_init_calib_complete(c2_init_calib_complete),
   `endif

   `ifdef USE_DDR4_C3
   .c3_ddr4_app_correct_en_i(c3_ddr4_app_correct_en_i),
   .c3_ddr4_ecc_err_addr(c3_ddr4_ecc_err_addr),
   .c3_ddr4_ecc_single(c3_ddr4_ecc_single),
   .c3_ddr4_ecc_multiple(c3_ddr4_ecc_multiple),

   .c3_ddr4_app_addr(c3_ddr4_app_addr),
   .c3_ddr4_app_cmd(c3_ddr4_app_cmd),
   .c3_ddr4_app_en(c3_ddr4_app_en),
   .c3_ddr4_app_hi_pri(c3_ddr4_app_hi_pri),
   .c3_ddr4_app_wdf_data(c3_ddr4_app_wdf_data),
   .c3_ddr4_app_wdf_end(c3_ddr4_app_wdf_end),
   .c3_ddr4_app_wdf_mask(c3_ddr4_app_wdf_mask),
   .c3_ddr4_app_wdf_wren(c3_ddr4_app_wdf_wren),
   .c3_ddr4_app_rd_data(c3_ddr4_app_rd_data),
   .c3_ddr4_app_rd_data_end(c3_ddr4_app_rd_data_end),
   .c3_ddr4_app_rd_data_valid(c3_ddr4_app_rd_data_valid),
   .c3_ddr4_app_rdy(c3_ddr4_app_rdy),
   .c3_ddr4_app_wdf_rdy(c3_ddr4_app_wdf_rdy),
   .c3_dbg_clk(c3_dbg_clk),
   .c3_dbg_bus(c3_dbg_bus),
   .c3_ddr4_ui_clk(c3_ddr4_ui_clk),
   .c3_ddr4_ui_clk_sync_rst(c3_ddr4_ui_clk_sync_rst),
   .c3_init_calib_complete(c3_init_calib_complete),
   `endif
