`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
OyK3b/zF6wevNnCs2nV5ob39gNM4l6x0djCu5vW99kx+sFqraWOzs9s6b+GrKJWCEYFkIfZK8A3m
qzwU8e5TJw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DuN+wcOZSyf4ZrkQlgz+YUYGi0YobPUWWEtOLKAQhWElDaayqNjhexObA264ACXZbaxzIRWhFt7a
Ix+3I8g9ok48gl4vstX5RoHhxpqaBFzOSExVPFXJFnJAxOne3WFJ8UOjtJXGOXpiM+qdnLtcG888
JfoJgOWGOEdY0/PNG7o=

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FgRaRjgRHYpy1dj3OP5irvjBcVTbof/xM/3iNjBNashYgSGBmMksFmXULzyxeJ2kRxZ7DSNDD9EH
3afrcLzsyy9NqEGI5629apUYeUtAma1mTa6/igh6BqU1nPJ0boD3CEi0uu2Y24sjRu3T/yJkk/li
g6dNpL8c7T6H9Air3PA=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
slrkxLi0zi2ofmPLJdmO89CFR1hollkJ+IUBa/Or8hc4Yk8dwu21Zu4fYKVK/ZZ5VqdcHN84TCox
muUQj/gwiwgRldXW/pLeXEEdFIWPDfNJXzPu/KRDWmKc7vgsi5f1YR0J6IfxQyaXBI+P4M6iDfbP
lWQFlJuMAPZZgCye9gjPTgS0DbJOrThk2W6mFoIMjPfgsoMEr7yYcdixUdBhiu4vc2HqjN0foipW
cGn9lpk587fX46BdSunckoRI1YxozMIu/y2lVyFjZXGfXasIyL50O4dNr7yf9fpIKgm23A5mLMOv
CW9UI/m2RwkHP6AHhicve1UjsX5H1kGcpaoSIw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b8gGtSQ5336bWU97rPov7OzSmu7oe/V0Yqrxm2GJJY7u74x1squJKWxTHExQze2GAmo0wjwmE4o+
VQmeWyDSRp49AgcBR85sLrXiwJIdrBWVzDMT8euM4gc/sMOlVNzXewuHqW3Q7t4HXJg5pbn0tnB1
9hhpB5Mfo9senobUX8SIdfi5fkWBlBiSArenQYBCW5OKC2/ZrCwJSze3h1TY/jFWQEXciZX6aFmV
AhyADOSWhlH9UYf5/lavjsxDBdSJ4ItgFuCIaWRfMrlXNSxZPgRcC0yuJVURNidTJXYlXoX2o189
cgCz2raSJMPwEAVmetrvCXvMw7yCcthmsikZ/g==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kCQ4y79zq4ueHhzPTTez6WplAFRL3JjR8EDeUZqdq1W8P2vCukU1Ill16jdF93f7sLd8e8bRS4/n
qwtc1Zzrt2+/AME6S695QImJiBpa06eg8qE1Htxn+aoBTQrT1PSV/nypS0hMdODDInvLch1jneTU
9TDCYXrxSLppHRlBaERKjji3JHcd6AykfhwZ7UeAgZXyIhujFqBCgOCW2X34Uz62B3eqGzi7CXiQ
zayNxn22i5EOGZ1D4kN9Nau/o2G3bIJep/c7sDlMXToUEyBpGl3kpDrp+sbIpyDA2qwNP5zerBzA
0cx0NW1Qe81yPkFYBVpd2Jel+ywwo/Lk9WcyCQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15104)
`pragma protect data_block
YA9iZEYrgtlhaFpfx3yCyf+dyL9EkFVIOJEcicWV10GGZt98MJS90OpQ104tihsktaJWbtK6nbhc
T7JNSdlM6ApMu0dXiEYl3Hn3zpaELMhA1N8IieXt/hqGwcw4mZ47LMfHHvzfqzhtIUXQzkoXKRaI
h2HRdaZRWpmxzzRJOvU/KkLTvo/VfgaFKMc0hcn0maNrThhxOHAKGu+fS0p/WvnluGwimsT8cpOk
49R+m3yzHLJgPSpD1fG+7tsFCvs6NW2m2TFOpWNKB0xC+xhiEJS074i2QTPl++CLSS8Y+NhPKABO
roOpHnvCaq9PXdFKzXt0NoNPYcRkaFgVxpOqEKm8s74kTbOTbgotODMkqtDWCyhkFWJypQvgszmL
AiWHhkeDwt1m6WyRGU7Gf+5jWaPXBMWGphewERzaM9PlVPL0xtgtqz2iEPHHMNoxOqteG7Ae1iCi
vUD7RIyOg9gWqol+T0f6BnNiKZYoa8iqVPoYF5YdGRR3J+iTAxBpSx4xQdkgrZf3lrCxZQaJDjMa
yqzrkmlEBLrNhx4HeGxVJbb4VM7Q06vJeKBVYCPumZw9OIKJwy2FikAs2aE36TI/eptNjM9ebj3j
CnMHA9iZinc+nlqQFqbJV/L89vexloB8wlZteNcQamW9EgIbUqFZ5jzNVZ0D4/1bo8r68kh8evHp
bhqMcy100jccmGh8qTH1TELslwUl/6G1y4wGYY8+ulymTcIIInSt+HxVitiJfaVSyJsskKRTDsUr
rU4hSzcEsiReH4W5Tut9u2VR+T+TJ2MhZmQCATfbn9JTm9klyP1OUNByHAILQohaSMlio7aoynDl
0ZUr1lA1yxN2U+wYRssTHEdhdRBmIxgNmKF1zeK/2tIgQmV4KKdgbqAFTaYLWjUf724gf0fjjV4k
DEyDbjIL2o1SUlIi1HUJCMswdBgKzVX4qBqlgOsyLSeD2zJGxmiI0DE4uSp5voDqjfepZQT1vkrl
bSmEyt5V5yYC0g57nx7K+DXv4lIMaGOhoiVJBBbJMPpc1LTedc94Uu2Dby1rjLOrlNScu6eMJ55F
JFaFq1eJxkoQn0189YqmEEJUB79xwg8El7s5sDH8sgld/VlfDMuzq8OfojUu1eBGcUnf+a8ji7Lc
zgG3nbViBhcY1NmvJ2DToW83S++KEarwRABiYuUgEOUDij5+UU6baM0xM6FNu0F5Y73SArBpyfwi
ZcGAKK0vc8g42nAgNPUNiF+bZr86ZTZ2HKd0G/Sbwzqsn4iXww58LyZ//34iO16x9rVjpIRzPYce
rY0njN2PlYtGvpapiA553IYFM17u+R0QrZg+Qlv38vgCITEcQ9P+jLIG4N7vfSDkTx+7T6/TzvgP
tomWbsO3gN2hHAWpMb4YcB07oP1i4WWQH55NIRNvVLoQw7Pf7CbYEqlM4CpuvjCyikdaPHwShIaE
pRh399e244LPi7YpKLoeOn2S9w97vxmiYH4FXiLhvbefLSaU8RYa2CBIG9VfT845iqoQI39B5VzH
SFkelUdbfykqbV8AhjR0/SRbVU9xcn+W1Aq8xf7ZVf+KHOie0+LGh3tT+XB1aIrVlE1Vs+pfTk9F
deYnPhdLTfXdSJ/Uw2T3uXLpuuJ2qIfzF0mL7C7tJz88p5oqeyahR5C3hsljDweEfA9ad9B9ZXzR
axfNoORzAwF2YBPWG6593IKU1HyMsSuGmG5cTAZnNiHbWEMqgAoiUKLFgZgBwdli7AP18OmSwP+y
LLJjmwjEbS1p+1qontj6NO+5vWPlJMIo4+GAVTVTDbVk7ri+f9LJcO43hJs4iTq8xXNPfZLctYSh
/Ras9DnpiNkY0cnd5hs8L8RvP0vIZe6tNhMBjYwXtp9LkwNCK+bpHnM5+7bKMlZ1aoxsqcHlMlRj
+gL3JtMraA7ROR4WqOaVQUpztP03QYq0eNnFkr7WPZvnjE8+nJGVwY4Wm1FQQHOOol4ebDo30sql
4kEWfsJlIax3w+U3JyPhjcUyeB801z2k9+Y6GbaPrGbjjAUSaRi4FpGxKRviQE8Nk3uGpzYsNz42
TnWtwrbM4WyEMyYxgeQv56B1j77ZPp1Vx0zlqTI9fb0Nf+oiiQGgf5SXSj9bNosRbf46XQVrx//h
CtzE7IYMAriiP4e7koLEnT5aTdIPWdV/1ydSLATOB4vIfBLmfsJQdBpXFMEqSlYUjUrT1FzETwAk
BaP/VY4q4ZviINvI2zWmcvxarNogXGghg61q94w/c0Var5lkFVHOvWUBU6XpTCcy6k93CVCS0jCS
Yi4owkNKbdtb5s8SZIuni/Lr6jDBeuT+14YHrf0UvuNmEGmUNAWOKeBqJK8sV4j/U8/RWzKwm1Yu
OZHFPa/xh/CZtR8TCzfZZhznfjhRzXE/pHElMFpPW0NJUOpParByx/vDEe2lPC4XZr1nBrQg/De2
Avwwq485VfDz4SZ78ghwN0u6w10J9kgqTOz4Z+IhxHdxqZ9vTJdrCF12pRngDWr74RMkUWYNG7gQ
O8R/6kDvPx3IM5vp96dLDtrF03vD4g2tfE2Uk+Czml16P/1dGged8yZd2Z6lsR7MP6hIgEXzaTNI
lnDk84bes4oFwAOu5YOCUdi702pE8Ncl+pqHTaojGUZPQJC378Dk0iDj/4C+FMWYX1c+A3f8jVyH
Y+5wKhCUsQ6fjxRsZAF2QmWwqkrmkErAcpNYfPsWjB+q6Pd4rlZckbpcD90VKQ88jwO/7t58QBhT
5lAAh0VPvXW3d+sgHoTAYhFUNz54oT6a2MjdkPyEkkbBOpwZDoCqw3xiqtdBUMmFHu3JLBnxmJgR
SDV55HlSHkfRGyy0jCjXyLnhS7TXAAQ1EiRvszRKfa4IpOL5I04e8idMZ084VzuQovATAlYN8J9J
FNHCGAV7uKkZgPeIJj9DKMhpRjOgPEyjzOdzf0ZASONSnqb3bjrxtpQb1ORloEYTP83fe8Y3FBLI
Mv3pNK4N9JVks3/r5X67G7DDig+hcZLHdiRIOEjnEjQj5q6sFj7w2cCS33SgufhojRmPCF6sWNNw
32TP0YkgFoDS6lUtxNKEJH9kOxEjSVaCJRfvc2Qp7bIOmRRWAGnYTkjVO2biayvNSN/L7KayccyK
bjdvo+kaYrMlSkK8ZPHDgROHIBud0ag3NUq6z0dWvifoE8omSkeRABuL0U7b1UfOUrzLxqSjdlqp
INmjD2g1IA5103Lkvc/WOkGLhzRI8TCTdj53AfL7PBY73lsSYqiMMbZ4UVvlu9MAOCqAemUHlkqx
NyN3EuQC0QF/Zo1Iedej0dSM/oBlrk3W/FZhg72k6bFUoyxOTqduKT1nawH5XmMTiBaDngJaPnz3
Ovwz26z+xKNB7AfXNJ5X9YBnn/kfnGLd4nvZ2010fRoePvAsHELRK/0T7x2/PJZL+GYGTKItcBgN
8mmEFph2C60OMAd0TGOFbupDLurb/GuhYYoJrDB2UUbEbOgZrJO76co74JO9dvJyInLJTOyIsI9z
0NGMxzT8lv5xwPpjykXFwWshgY83UOWLWhW4Ay/sD37zlhZPZbqOY92ybeOWINY4UNJ+YjaB9Uad
jlcmYE94sHf8hEAK1HEDZDQznllAiCx47hZDYKxozkaYeA2Tqa25QuqMYQUlInA8QM07HxFjcwzu
6XqSHHxNTQmN29RB5cN6kflmOAOcVUIsIlchdORSV8H2KOiJ5JtUdxHOnbp/H9/n+u1JL+i4USTP
witaCRsez554n2BVekT0KssIaB4uyo73vXMaEP2MgPoXbij8p/0Zfxrf84UhnCQHf3nn/o33WbaX
TMAglw8tojIQ32yjVlmTZONk7qkBDZgjSWFBfL/ShUkZ1c/TFWwiR3qRQwzz7Gp5eB146vO2VKK6
zr+ENwbxjXqudUesM9fuGfauDuYPih2H2U8LX1mrfP4KLL6cPfZnfPwim9HBfx1sxncFPc3ddqDz
CcXehrRH+8KcqhIqAEjVUzlbsz13AFDBoUJnZA00L5JAxRauuuHaurCOahqgLhJHmTvIbbR2Wx75
5O//1rjmy2DLkQ06+CX+aHSEarLW/ocT7aOom64fMK3cerxkyP2dDg8VHtbp6LyccZDrOqIAOWTg
k3ddvvcKX2c7rGtKt2sWo1ClyAqELhtETQodrV08SLciIiDdNexwXmc74ZkdBRk9B29rPVATLlCu
0/gEh6gscGKtHUQmhQssEOReUCiwgiBI5NLO/lfkraH8RKdodsxof1eao9qH4NQnSUtKJttQXdPM
pMBWuulL6L3QLPQMBlAQCklA8ipHzc7MCoLxKAYQV6n3cn+M1iihh1LuZ4+88lwdaotvom9Ee/Q6
QmNkjhcER/z2eOVLEjtMiRQajgiiUEOOchoQK9in93LTICYIKKEwh625unubbbxd3pZJzeD7bxY+
aEO5N/1LkKEFO66VoXd1myfdAx2M0BXQT4TXsLSRMQXzepT0lnE2Ji5RgZr1fCPJ5wiYXUPEWH1t
7XOhrHrokom5gXQ5Ah+rewcl3fPsGw6I4IdandaoRcVvmvAZX0FVx513U5jbYckPQUYmYPYLL7ZR
Lk+uR4jMY8/i76UHGDaG+NF1FoJrOu3vtcGhCkpmk8bt9MNI3eKNK/X2JF7Ndl7YrNzVrq0f4DdM
/oS5ENwDjpHxXCM19zBJ47bXUcWFQ/LxUjGaSSzhafVaQcoemTsR5EQyOrFrxhcvDIUKo1oW79k4
ohZdgXtPsja001dAAPsBC4C2i6tHCMKU52k5PU0PzCfJmNM2acqhW5fm3j4sJgqqbLrxiIqhBttL
P9Diyp1M7IaAKUrQw9vFmPzsXzoVttMGr2hOAjACqWgbKQt2OuXiiegiGlwppe1x9hOkX1QlZ0Og
0XKmpU6+oEvZMFHH98LbzKKqRMjJP9K3AMOfs8aQqwpA9nZtmq6uW+GBswk27VGhUof739tXZDoB
+BoFt2ZihlgoAWJ6mR0tS/TAcL66Xz1+nOHABQPrN5E9rkPL1mONHSqN7UD9a3RfnYnQGszQoArE
BZwa4/gAY41OjWVTXnGktnm764KCiOuwp5uhvn9N3a0dWcdQHb4ee06VxuYWNlKYLDRFqyfFcbvs
vtMoooz1LZqIogbKeFNZ8Sk2VlvJzripwZFtd1lvGELXUF6YZveRnFsYjEocd/MNMiR4MADN+0v1
yXaAqinR5QCywR7lKBAIr5WHRA1xPtwxP+8/8Qag5OvPLBUppmcCuVTRLssMBESM3SqpFczim2Uc
ZwZsD+UDcDR6tmDNMnUPcUWKUOJeA90i2Hm6VOC5wNaxgRlcswjHG2f1ygsX2lj2Or8gBKy7pxeu
0CrarFj4Nkn+zI8HDaLrMLFPeBevaH4cciqQkvdQ/LQJaSSEi6FnayQfzPeAVU0MesiUCxV83Aw2
I0jc3Uiq572oJkL/fJehy3OWXtyZRQ6jdKl/2BbUg9XE7u9iHa0nDnc1t+h+I8souvuAtA4wUIQ6
mvJx0ObWZtSU2uQbzWE6Qh6uFVYFBjoVFB81Awqsa3SRJrly9RKdRAqyGs/8GXiFqUg0TQtv+lJZ
UQx+8hRs06MocLtW8I448K754Av73zpbC8ijE/KvYzL80mCn5tmihUgc2U56JJ+DtZpkt98gl8+G
TplzU6326ighNm2KXBx5vvXTPQREYMbTfTnYnF3xYqOoCyDUd+Ko8OWZomO8hxdFcyByA4I8Mj7C
ne8RiNQgWopy8wQYTJoQo2Low6wQwrlGWW7hcinU85ybqG59a0c8pHqjfbJ1Oo5MSUSArqHwPKv1
LQE5EGRYWBHRjk8ecLc68OahroX8xIJ1VU2iHkI+T0/YthrVkPbNcV27rZOpx5UM6rnSDtYwHwFS
VOa/x0KLbp6iwk/eDLroRf+o6XVqvqc4PZv3/1JDJIqyW3fyzYMxVg8uVA9PoRWO8TYGIWTFW6YX
tZWkd5iTSrMByfsoZfAWnMcowICR9UPZLlvXZV6XP66Mdd002oPEnAueiziPjAYohJ7HlC3rft83
9RzsdKJkTldZje7OCcV3jIz2y3TDjcOqOsbayRwT5GHLeaNJLYqMzdWJ5STPH75eHySwWHFYLGH6
R5A8ynEcedfI5PN6Ubu5wrTIn22hGn1fyRshvWKYdePItemVF+MGZxTZ88tMsAmsP3Ee8T4S89sR
83X9n9bGb4harl+2uzfy2MxZZEBhidq61pkAjMD57w1sccet3DZKhadlVI+ZPwrRSHXUgEIWTU9Y
5jhei4qlrdyRFsVX0oXhKLj+3b+vypIloYMb2Eq6wWrnYon7P7t2syFfGnoT6opTVWuD9/HlnFAF
/vc6P1RLYu3w6KqQUk17KimcPi3kkQSpjiYOkfL/fhsH7uu4gmC9MrDZQQnsflpdo9BOe/+O4nJi
oXg1H0Yik3fmAh3inYyvbgKQhMrQP1Wy4H3EJdeFBMnmc4afbyjzy3peq+K8TduTXnuFlzrWxvPD
Jm9daMG326pFXpWiLCAUZeXnSE5C4hW8v3emFM+VNlM69sWyob+3JbQ56QKUF+94p6cWtlp21jAf
B3vrEBJbyu1sr7LPJbRSIBFu1rQw7pvHy7caNsEszHpItMQBL/n74Wy9kk7dGc3oB7xuY7pH2twZ
paUqxWNht4Lr0qRrA6S2or3FFwNONOLJ7rP69w0SG1YE13BpJ2XEGpmnCmBhz25TG+meXHeFnfUR
VqaPI6m1Y9oi2FFGsqFLus7+alKNVl0stuAVQ6lWLmHBriJ3YPkqvB00ZUcTS6FrkfYp71jG9iQ1
dW0oHDQbN+PLXEAFSce4FelbZ1AAYjzq6pBx/WO2DVGE9KAIf90FA7zfzKVM1eUqA8pWfLNGltUH
XdFhM0NStA3As1N0W4eQnMjiv80LXkazoNzTMycl331StCe3qOdH4WRLrCZnU2j7hrLs2yC5cbik
epmeqRJBSQ4mHyiE6rOiacqTlYG1toODK/2SB3qLjevlVKq9Mwojgpk1W4pm6Rvjv0IUtv9bdw+2
ttEng2s7bJj6iGCgCGEZocfOBnr1RtKF4fhIGc6SeQMp2+JYXkzTRUC+uVlgi6D29/cIROAUEoYS
NJ/bM+IPZFi18qpvek/m3uUmIdeWmX/cxR2BZ/ukJ/BsVjGbMIPIDaubMDNKx4PB6YdZ3okelzsz
ysYVbi0rj+EZGiQPTxLabUu5JKa2p8g9YK8zKjEgmh1mY3VRrweF4nrD3/9Zn/VpL5tpSxfoqvlS
sTVB1NOoOsjxP3YdR/ssb5RPR/3WR01N2TDfVPk6seIHzg+8olBPI+KXr1rnSJxINvbCvmNxk6vi
VN+5D4Ah5qO/wBYhQZPBcJKdKUpbRRwYH3e6orPvh4dMTqQHnOSo1f9TJetaoc2wPuJTM6B/2UuD
AO+g18XrXMMnFPksEwC5UyGDDtIlhRuiAhrMtCaxGS+z0uWvryGwz09WvUmpHi51CfhWf4JA2U/C
OZNp0eDTRKHH+hMPZr8xvHB9ZlGuQ/epwO6Ao96Xcu8V0uoRtd2Gbj55AIQytXaXmO+PLHQ5UnMs
cfgHnXjmklFgU7uaADwbSd2s1ae0WGlq8hmITQTR7clWLaXYnUYUego03+tDDGTqjuqUbnjW57aj
lrKhRSpbokHYZy9Cgh2zPxkPaJ+AbwrQUfWpLGStw3UTvZtWezdjTfG7b7iHaNXdqGsPDUNK3eqs
TpdWEizr/+cGNT47wAH4x+zbzyW0PcX5XJnxgrK2oqHllJQ72ChLbLk7Nf6GprVkFMM2Xu1tMi90
T5X6pfgbJciKrTa5LSWRvArwX4abrNrmUVh6RXBXOJJC8VdtlCpo7RvOwi+SazRccmtatloSyzqQ
p/mInO5BVKjavAOOXWYqayn4lmhj3cCdEsYuZTac0mlFvC4q2oYbv+nHkYOgmDCwln/xM0bZmMBF
M09wbw3AovErYaqtEzSkwwXZeFDgJtQ30SI4g2wv/1rUBYmsDxVBu/iZtOucSdx1AcKAKQoKn7Kj
nADny37UAhW/VhxjG4Ar/dNDrGh4o09kZAYxJsHkbnHFow157Jaa4qcNDud5Je3hLiIbNDGskHum
qkF6uGny4WNRDGJY64lX3FT/HBdtJUClDkXJOCTD1ckzUthOd1YUjBDiJ6//oXvvwhdLrAqrmL/6
YrF9sFPaOmJa4q8ssyfqarwbBYgzYlaB6qy4PvXaqDOwI8QK9HtDk02dTCVb0JT97yjyxkq1kWBO
kpN22XN+XjDbahx7CvZu6k9Yp0Ge9opwN/+5E/wyV82QLGuDEWkjqU+ZodIfZg3kh10cwQcFvyOA
1Rt33rsCZrmSEEE0aW4/7wghvaTHHLvP3sYNOXmpcW42dp7Wh+euvBodgiLbO30YuXrso7FUYq40
RK//zAGEyd5omTELp3zCpcsi/saRHSCSatAFIwZBQef6niRaqD/e+if41TrU1V4j04NMnGnO0UNu
xbYGlLQVe4NA0OOigTvT/64+StMc7nIQb/44CDJg4kq+b31WaFJNEo0iOwYj0DQGAMgWbsmDpvY8
bn3U6sFXsGMuTnUawHXNEEg5NsNd9lv6UHPEF6tAf4uQv5q+LzLQ9W6me7As21kZ1kNPoGMFIcl8
kyTtU7Vi0a5272HdqSDn6eGsdpd0f1J5DEDJpLbwpP3SUqGY8X44fWIxlxIAEhiA2VSc0jYpEbZ2
iCqoH1wgkqMQ0LXaR+DPmDSqq7gmQKlPq2Bzph+39Pa/JzXt/duVq3h15cdtzYcEeeYCQvpO8HUY
Qwff3uuoPIQNfb6YDgjMaWhnuTUpS7YYkxVC0xxgSWgOJ6HGqyrFHHTOHrlanhAKc3jpDLt45emU
G29nsVzP7qA8r5uR7/r8rcG1XHflxQQ9N24h+9SwAL3TF+IxyDa8yFzA92s2FTKL1Qn0OnDg256M
/tr2q6aN5Vq6IRJN/yHJ/mDsVDGfUYnDTYFw1iOd8kJxjUh3AkPAyJr+fAbvpDCptfi3nPQVUyLh
ClipkY/n6135NYrOQhDj+lAh3Jk4au9uCzUhYcyqmTYbhbeUh5tXc+K/f7N4kXDbZRHoyF8ihR3+
NcHrKxJ95y8yni/9fRx7nV0jnIYL06WnhxCsar+o4BzsmUVxIaunLUTf56BqQBtcYyHL04xQ5cCN
j9r3JjPmafNks7arr4Fl92FJskyLUBH9Jc8KBD8ACrX+2KeG5ACBDJdcjuHKmZCceKLZPRFExurr
BL6gUp/xypJWb37l1zc6n7qul6ciTNtu6k7ymlV4me6aKAXSCnDy9/28TKF+cieJ7SaSqGpa3CB7
DSIla8e4vqMlXxWz4TJKycEhH+/1TcbetlG0lVwfvoAeEiBO0HE/Pqx5uOU3TwLNxLE5skhCGtJG
LqhDx/miVByZnmBtTMtt8QW7V+9FEkD/stm4OcaJ/SeUyzOKaSK2UGenW35Ukh9BmmqZT904TfQn
/EzBHWpWycn+p5ug+HjgAyrWzM/tSMCCRBPiUgCGzE+HwqAXK8TprlAIVqINY7Ymsj3/MokReyqB
6Mc1Db6mx6Q+ZLevwY6yNecdM1y7vlTgVNgU0jNDwVbmYNSoj5wGTKxzU0ctGbtofYRRCGONkE0P
9Nd/LK00xCbKE5dLCiSHpINfgDNQeQLglcMXFXoGJHxOdcNVgICZhHfmotmZRHrgaTlqdJR+6koC
ZtAgHkTHr5uBwSAFRohlPQEqn7bq6hljp6d7fdgpyvJ2bwuQBcKLW+we5T6pzc42/fFQAY3VaXpe
jgKYq7hc02nQfOh4/uw75WAM4PmFAgQPLhPA++J6tGZYLtz1pXCO6vYNufzJCTmw/rndf7LEGlCQ
F9+IcsfV0+00yOAoRDRYAtb/kKfBcCEw3qMzBz5pcrvbWOmVgEX8BEX4kcCk11A9JH1ybY/v6YE5
02MO37h+N6Lq1No0GC2oJn9A95tvxLspHSO3sDc/x6vvIl5Bc1yEuq0r1bjyZ34KlxSST4zn+/vx
wRGjbLT/kSjCN3qwY0gyb4UPVgbDUEqJLZmpwixXUbicPYwtK6ve8P/aqXB2v1C8JOt7wzbXwRiE
hyf9mUBEw0Sycp3YFAZ4LqquPjvG3gMRhb1GrMNvWilODSiEBewinfajOmv1xIQUW0jcVTacpW++
Jlelg0rOqNPW4DRnWRcfai5EOd3QupqqKVMEWEZKFIrKExNewZjKQkHeS2qpUwdQYkm4mWRNCrdR
gECvUMK4wt5jdp4e1GScbixZr5oI4CEVS34Zr85/uPmYksBRB5xFMPIXW80mjOWoyh8EkNtbo68/
PW2XyEiE6+P8eSi0rzSKEbwTLCQt0GG3Ew85EGDnrlgIFnrrqE6E2d5Ei2sc13KMGInGLTByIMJd
dXsl0wdGQ00DpoSx4aqWEzgKiCUdz0QiSzda6bWSlCrGnu2sxy5fNxzwVSB0UMx0/B0Ix30M3+td
18C/rHHnHaDKbQIIyg54f+Tu+v0FKUOU8LItIfo+5FIRSkrXWtpQHzV+jzBwNDN5IPrykKV4ScKC
nJNFFmzjIdIwHJu1YyAPnxsNwdEoD0VBapslbQKSiWHid4pK8GnJBQmohFB6pbvSYTugqW+spKVY
6/9Ln/CANnEKwl1w7YhVvzW4R9clt3b3ZCVX4i2HxCMWadVUwDuduxx0S0kNJabIzAlV5QwmpROS
XSO6NZykgoYnEgh28sawCvE3wZMKDCIxREXvnxibUypp8CZtv5ae8iaXZkAv1Trixk4pcbdxDINN
03owT8xShJeRG2fWbwbufZ7XIJK4ggjIspf3dlidRccu0BjZ+2If0UcV79xztMYGeuYQoqLI9Tls
LiFz1X6ypTHQUQyTWwvwqWcltw1tsjLeZRrtCLWsYyXAFQUP54/EO3vejg+cr35csA6tUKL7+q7Q
lYUMwnoMgHhKsJYi/d0H6iQsR+HArSa0ENor6rnOdZwmLJKoGF4fMUFiZfHM7p/kXvdgXwEKxM4v
QSioVcGBsIE2uj3kQ9bDDHyrWsTlo5fxcMp6j95EeUvZw0uLvNSbqNphP/6m1lxTpriCvuGXR89L
x3mk06+G2stZdfHxgjihj55o+jTDHmb5Vsj0pcDvbMLHJAwVKo7FUDpwuLIRSFFeeNvzANnnb5Iu
r9TceAhhpfcUlE3pPLklA8ABhTKRNXM3qrXpKQGxK1McDlOquFTz7vDi75GFQdPFc4e2PkaLcw0t
F+1BE1yjy63wAi2+QmID54rfQTGt87AkawrhVoX3CZCr2NxpTzppO71BFGEeZeqDJMtL4mGBKfpI
Iz07v9MxwSprBhEFApTcqkzT8mTJ0LEfO1Wx/YVy8LkjmA6+1PDuegRHovdhsc/u5IMkTQg/HD1J
KBOlFbEJM0zIUBj1SNIgOpFjt0MlX5DP46IdRHiec/5/eiIyGYbns4mQBabXo3/DbjRknsGmHgUB
ibIQA7Krz47WBVKwIMJhvptfHr6kLG8CV6cRmWgu4gboAhknlvkhRiRQPC+dJaZmoa6njfcC32Xz
+6SisJMgVkI4UNvva/x8/yu2SnCn7/C5rf3KPX4dH+sv2uX2nPv1wEy7awLlqgHm36e5q7hrK/ux
6K1IZ2Yh0vbK1hZ3tKRBBm0xfasJAamavsD9GkRQySWOcQJ5fYVzYk96KqYgyxdUPQKecCanSwPL
nvDCCfNm0XZZ4cmGwgyJVLncwfa2v5k1eusyV97oEgYh7+fhAkdazAKvQsJVw4oXKDMm4qQkwa5f
hXzmm0aHc6dGgjTbSTXfgFIXTyD3dMOdaMj5ZuYW8LVR3Hhdq+bR80gixwteY1R9/+qMTqyJrqd9
qyNTHyfZpjzmhB65lGD7vcVju5ukow40FiFu5ufKmM4q6Kz1B1qccBphSPbjXy5W665XHqgPM0mV
SrXT5BztJzknni8Rtl2qi3jq7G+MgwV3+EeBnJUNmSBFlMAJrQH87sY3dZS+/rXw59UQersy99zs
tNYfV1f7KiCtVaBEYDsmQGb89twCqR0pnA+nVCOWt4fHXQJrByz0VyJsRKY6hh2f8m6H1ETwbEs3
WwQIQtU8smGfbxmUQupaGO6q2/I9Td5x5fVVKD7VuKXQGKukYRvNUtGpw80V7tldje2R1SFrS+Yo
yjf8p6GyvSZV87dHoCXL1gQ3ZobT5yy86HpUApMFK3AeJYh8ZL9qxWi7cb3s7aIiTR8PzNXHWGWW
US2DWf7GG7Comq8Pi3JBIKjGkahAgec8B10faYF0EssUhFin24TVMwBE2Wpc7J19hKQsqBJMPAYg
fkI/obHkM39IvZT/HL+0IaKpt22CXfLFhnFFwO9dDJ4dYq9DM8TUtMpbyWhRwQTq6OwPWOG+QvNq
xdxs7D5b6+RkxvdcmNKTibSXOr+hr/SdFcPbLlKpky6miuR8GLuo8Gp4rIiKSBfloRSH7E2brKIN
fZralVNouP92Xu+WPzE0VTtmRCL8ps1YcLYjwcPp5Du/AdDF3pfsDE89F1DrrffKOCsmGpGi+FyB
fuijEbQAbDvF8xtH4LvQJryDt3/nbQDkq93PG/kbQ9S1Sfvc3Ynl/vPHHZXZ0DhR6mdb/nuzwW/U
n54hhAViPZlS5QaW19AVCRINC1Ws8Ifsz0KWxzF+nHNbDUKeFTPi9Oe6ySRVWQcHtktea5TwmLTy
Q1nfKC3IP31J4CN2rHIxcrSeXZLxmZxMsk6/hE8Va9PSG/dOZGI/eBT39GhuxQIdpGOmsZnj2eqA
ERqCt+YCrz3NVCo8pw/cRaxhQIrqtLO4PkYPhJ6szYUu0KJj5aLLmGk1ZP9LlrJ0V474cbOao1oH
4IYMLo1mKsNBYXyYF0aUPSmstqprHX7kyy03yPj5oXCi1RG+YH9ioW+Rqi6zAYkqwMYJNllKTbET
gZmZBaXqB3RcycXRx8gn8Tl3t0vdPPldsKylijBUmskCnr2XrbNzQVPpZBAGpE9azUBERWncczES
ks5nlIdfnsApEMQ/dBSdqvMTpcK7jD5vB5dCrSiTqdTnuGT1MCCZTnqDmAr9Ml/3VF+cD4ZJAOpt
G0ZMmCUqu5LuXIUJQm3ekVLG/awzisIdPs71dl5ZDGrfirRyYlWdyVeb93L01yMicbDBiEHige4Z
WLFdiNIf2IrqMWoZYJPA8XbwU58VUPn1TuZr1Y3qbayPCjx5xSj0xOcQ273pUuyGXqI0Gps9GSVo
iyHknsnaN4i3qKUb9kAp5t/2VApKtZPaU3onm/Lky5EFrO+Guzmupa0zUu400TfVGrtgww5B6DLm
KhkKDrBV2jaXi2vybdasPGSpl8MM3HaVSokf+lf8a+T9fuFwyztZot+KiogceEfHXJewvpZvaY2F
MW0EH46sp9tbKiO1KrVPR/rKsWGRJb9nZhyaZyKWsUqhzVbZxafI7Nvw1QTaPHIat6IcYvKTF6+e
ehIUCyePZMjlfWmjK8F+Km0xy7wgutjUcq4M1zbNkeOmkXkAzk2e/cM1PBpuriEwCL0OPgbKiohx
oa2aGtyh/RzPIqWr8jMBvjeGUo6pmaR9fDRtO6Ly3cvkiGDyezieABzzO/F1f8Ne700Od2dofj2A
6O2Lp4OmyPgdoht+Tut2fnGHmdCMg74KGdsPVFzwp8fWK5kkoZ8ZuWQYgsHvZ04Cc0E2CkM9ytk4
QnnVAWcZ+Gb7D3XQ5JzT2eWHvcSby0ufDZDzvGxqcQP2tTA1zEbe/W3mVmr85nVU4/WmToHK203Z
t+PgQ+u/uEqLR946svnwItRxNA16NhvrM3ElHhIjqzADrPuXy/d1m1GhKWT4PAXKHK0pZnnaKTXd
YyJBJMnE/bx3RbWkhqpr5fyi7VYmQDjFbq9AJdzuDxNfY3Bm0lOpo9FeRsYMPT6LJSZLmAy6yVjW
v1+BsVNJsnAzR0JcjubtGLfU7EVFCX5xkwRt7xCz0/o2Zwhs8w787LBpVE+4cJf2DSlUhHGOC/Lf
1wteMOlrICQxgCdgfNZlfDNHkbJrKeWFLneOVVYBEHaOmtkx+EH8i247AZcp3dzitjY/BBSghni/
/L0Z0umvNZEIPvKJiLPa4hq62W7Qwq7YZNOhVjqugNa11EiATWVudRjDz+3+qfkzckSBirD0oDOX
SX4HlfZOUEA3/GSZ7uYmotN4WRmevy8B+tqxI+CUfadLnk1+b70z1fY1LTb7vO99x5gdO1b4JOWI
qMswNUKHJWvMRS1Nuvvuzb/Z+cJ99yhyipFNJu8RBT9q4Lm1OxZ1gzX8GtpOQ9em7MpiHq8GIa4s
CkwcWjIrAyv2tVHGdcVvGoXId8q5D+RTdrpIUN5VkrwZSn6GN8g46gT8WF/0tNvvuWk3vyTZSP2C
AP6jtx3Dh6+T+XswHKaScPuat8uHyK0Krt8kBJJeGfUzLv9QEz7IWjQR0iKshCYpY1HFpv9yFDJC
p2dDyFQQ+qm2DQJ5LJEyyz45vCwcYrXKV+ybW7ZVALI+hpykAOCJX5DOHl4XXPMNgVNEsyfy08ZB
vvZWBW1BPs8q+JIOqH715oQSW8HKAzaAfvUcwAQdswHp0+oEQbs8WHWD2cHae6xRCA8+tHD/tW69
R5vXEGPlrn6xEmR4LOX62wzxOeeiRtpjaVXYxdoUo1P+/gkLmNDE4nKRL3X73pCKuBAZyS3+qLTZ
YheAwA5ljWcAUFNcwn6Cut/PpTZgaIowvVeXVH604IW4vsUK/KcXAaGTHQqJYnihcSu4uizo+sFH
LZYibueHGloKplQID0HJrJtjLI80D4bHsQnRcmTc2uBnWcRdUdw7YcQRwkafSrUK748Z9hXgytfq
JryDwjFAAkl3JOxfS5nEPrfWYTP/w98c15knUjAc68232VIqxA2qb+wAcZO6FC8ETFkL5st83a02
nqN8QcTsF/41WUy3YXEzeDr1c4o/mdcYSgZ/o/sx3+MSzkBfqPISYViE3Y5SC6rEjuwttPHenraX
HUes0zSj7j2z7l/XvxZYFVrCFssxT0hem5EI8a3fAklzWYnFcw6Zq1nyFFnicRr43wedJPeIgKnm
pTQklSvQ98iqvJXqqtq0ZV7oVhIeWpfTdsVJ2VMeeKiaBH20W7RgzrIKT/zZKIh3wXqdT1JdR3kk
PaVw0gr6hTQIriMT6+cVrXtEiGGwqP1FNTMiOYnl8WKdcgeP30w4cbKD8MuOTALljpHeAS94K8Ng
TpQN9a44NMWEV6MRA9N3Jjtz4zoIjDRTIrGR/e0IEbzFbt7N5Au1cZJxb1MWyGRjcQQpAVTGbIgb
euBq8lsBLNdA17V94DIqe0BnIL9vu4levG0g7ZozdD1+a3F1SLnbwGecuYs5mP5Li0c6dt0+ZxbR
GEyhP2UofKTxgPQ7+i9hIa0QHoZwxs93XkMzD9iahK7NHumm2pafgVwLqmtGO/YCr7m34K2yYHh2
B2Fuge3HOCIewSarC4qrxdt06sWd9yU+NwGa5+sB5irxIlV1qcQLKeYzK1D7Ll1fcSdT4Zw+I7ul
BCmOjh3HHdH0lcXtnvK7ua4UZ9PVDTdlRM38CeTIaUyU1j5FugEPj3tU8vmMX8Ialu9Gvt5aLd37
ct8z4c/VUnK4Q44rIItfxSrHRBA1T18DEJvjMuA9a4T/YDOfj1L3DVB9ENgUpPTTZOV4WYwq7VVY
I3TP8GSqKwhpvtZ3yaY8E+fUT89MwqtjqotiWV2/vXU8Oap8qYZGwgKaeK3T/qdixXkXM0cQcjJO
YEW6kLhfCFW8Un0HWc5NTUT0vypL0dvzblCDbmABldvFb186kU3Pfz0lDV2wMlXYjGNNx0GPN+HL
5VEez0vPn/UyZ1Fj6AaC6UwVOYjzAshgB7Nu2svbX4ln8dhGMyfaKql6si6HEc++1/cLIDDxBM83
L8BuKWPlZYiLrJZL4QvGZedlVb3zGils6SJL+mRnnqnM9B94cGudLugtyckeaXRtk+kDwYkayuRj
2btSLCKGUDU3WoTZTvPQyxYTO5e3e8HwxvTpBIhK+egMJIllsmyvjQ+GiKXUFR+NMHpbyQaOh0iE
0AYtDCUiQoXCOIUTVivTOn0QjWNJtIviQA+oMYJz2nKHduD5X0sIBw2G27c1TQxkOPAtn1W4NbDd
oTbnPL8P6wESp6RJSVWbITl/PujsHZsNP9eEcehj7srBc9pcYyLTBm8hG4eYOrUDGNxoP8V2nwlJ
joboy3JUItH/lqsBGQyj9eILw5r6peqD6OA5NU4zRQ7QNhbOYKlJ4GN1MhlB39PyzoObRZUR2848
182DIOR4PFdGEnI1SDP6AJpnmRRJxNBbe6AKjguZhUPYpbExidL6bnYkzy+LF5sKnfUVrBkphWRK
vrGAQKZT9MZgPrOWaLjL97pkn4EpoXBtLkPysS3GfS/zGK1+jp9cadFD4T0S5xp0tVY9xqPY5Ng/
KxeOFHvVTLB6ms6vFv0WIG5wVtJwFr2pEQ7VpWxozV0i0dB/Mg9z5kMipzAGsmzqs/3RVukpQjcB
9DHWqLEWyYtdBs1QDtcWlJAGQMyi5QPyEq1HLwwq2egjhqJqSbNzQwfJHgvTsgzSj3IBh7/AnOIV
33W1TqKu9z7xjGYV0ExuJUEP1DuD1JfqAqkFOR0ndLSERfvMaMPMUKki6jhkyObK9hkxTGYjsvca
I3onwCFeuiaj6jzGXNvQkPXDppKI9BbyHt+I6BwonOyx4IQfeyE/Oy52nuAwTZw1VR60xkgXZneY
+07heStSbhfWMDmDpTgNLAbeHAEKL6NruNIHZG+L8D0LpgqfCwQu0ObwIPsx+5LmI6ZNAKzYVctG
J3HpH3Z1rL4hs62xZoa+4OATokRTCpNC9aiD5RbYG+PvxV3NlBTQ6MFfQelsttj+/cr5jGzsOkBf
IPX29WigSdoEHZDuZtStFIadrAcQLwAibBh8IY/oHWr88uAXXzcCzsq0wlprPlhQ38dJJstC7c28
pO+HvAFCH6XRQ2NVK+mmi2mMd3ZIP1DBGBirnAzM0MgUJh4ulEO6/gNsAbjGDzeYOCQbQZ/sHR2f
LVTBPWJPhiFRLlqUJIkYxfjTP+Yb+zBvpNcrJxQRp2Dqsd9ghXfXY7D/vzPtWd01hOZETIOpUViY
KksMdMCh/zEudQ3JnvWNIk1BK4ujSECxCm/GMlK8zve4L0v/HgHIG8dGn3M6nn/b22d1dYBFz4mA
cMQ7445HVf1tthQOAXLPE0HcGCP99wGGk+i12JCIJ8N/ONRGh7kXQvi+T0GR4bBGHx9zdGT99FIl
Ioo6HnG2IPKbI7NW3rRKA/JSKsJ/wM3TkFriIPUoO911JzTzS/1TJ8SXHCoY2Y/6HJiKSZdJGIKZ
trEUZ8xBzBTsATn+AomswikzWJNLQ+nfVd/9zSyld+6coZPox0Xnm378AdOcicS99TfjjdVhrcLP
nBLlrypv5/+QyC08vCCcXDBJJHK0hrY6MyqlAYQRImj881cRqlx6aWMJr4J7jppw4R+TZRZxIGZD
o0+YCLxLo/Ca7R7vX0zwpCSZBPKQ30JSPhp80EAvQn8RCEMZR2A8dYRyYjqdU+cIdzSfA5EP5pul
9LhaTRY8DhyWZTPTlo93yiK+giCu7O7bMQr0kyWRprmOIaofFGZYZAYvgl0+g38nNLRcoJZkT3q/
amDu4AoMGey5cXEj6jI1ZWgrzbiOXKBqiMDWIJMcTNppEuny5Pch4u+DOsqYBZTkWoSG+d6YjmA6
h0jdNB0HPuHSwIf6vxkQWxTOGmroa8EjPc+dUoohSv7YHMCA2i+2EK0u4AZfD8UFaKPzllznrnP0
2JhHxHZ+F3zhkct3R+Q642RRbjbgkgni4vhQ8R32tb/wVj7Lv8PtTY8jQTi5T+0X7kw9EKHdSEgc
yqui/LzDkS7LN5l6L2FfgKhga0J+GpvPSYMoUzZMl6Z1rLiEDFM+7V8CAm4YGxr6VgGVYgEyU1NI
eYH0zyCxJ4YEgSfR3l0iGgXVmtv09U6qmMohX6BCQ6eV8n551rHexw3VCCcnBKZbW6Rs8kz5KPaf
decL2EwZJ6ztY4tOf2xeyUbZ/5eK5rNRAr7vrIhvE5UGvKVHUwGRlsZBVq5WzjgyL/N0TadEFRUu
N85DbNUCzhiO28Gq/sRTad4O3mHL7ro5ItACkA7MRLJ5/QA8THTo335PDinVK/JH8W8f5PEILvL1
bJRKuHjJoJPrbaLqlZ3OUASdwIxEtdWkoW7uwQcvsR78F83JoVCiZlmxLuxPqDps7DWGmloa5Que
3ug+YE5JTCcxDk7qR5C6qfNUDCA+BvgJuYPOGoLEH9FfOVQmdUnfY0MV6kbHirBXF5B2icNSt62k
A8e7o53x1z0FZjojtRZK7MYsF5z4SUhs3yfjnALr3zlfEHHMLlV4O/VfEWsWV0OzS9yUWtrZzomS
W3nvZ5nhhbEWxXtmqCY9rN5Eji3F69IDSrxriGpiCMkcSY+spj9jMU7OvwGaSlhDw7fNmPnYvkEo
b1Vx44xDMODMVbz4RII7sXOg6xop1Qka5D+c8uioiLgY2Z+32rEam5OLtIkGzeQh3cbqUQkN+hKm
1Tp5GPjzoW8NBGWhIMLY6/tpgpOogFhbibKUNunjlrZgtV7jhjs73zb7U9jb5EByQfQqqRWywJ2L
X/jQqNDZsHGDP/yDLGdFP+EQNZO+c01TYanv4HVxQ8e2A6w6AS8Po+eaIJrpT3u45y1xEDChR1VP
thXkrx0LiacfnVTqdrHFPTXxLx0M9prQFykKW9n4uqZNgPZFFEO7kMyfuu8saHAbt1HHnXvUff3j
6Oi48+bb6yZWwXhqF7nJVxML3UahzhQZOMLEVta7S0uHmlmsOYkQ1GQFoouP8aQeTGTMBLwffFOf
CKeaHmebz3AA3ORgXvQ3Bb8HLPAvihlN3J4A4lQx/U8hAEEao7TevFcHPlDV3DFC82UlEEH5Vsbx
vSwxlxDMBPKqvBtArQU4pk2vvEh18nP4p6lw3S8FtbSCklDy6fUlLlaHrp8MqT07wc/e9O/qKrTQ
fQ+QxFseAv2nm1xemFYQ22abKcb64cgxmlKv+rHMJOqcktvaH5kCURTsXrOhg/qC4p8rgYiHiNNe
mOcoS4Gwm5U982Rf6Tzo3IlP91l5HgogtGT9brTou+8+UEs4UFzUY7q6MXeYYepGgscqqBBQz0Z7
wfp4qW6M7jX7i67IkRGzKJt3oIiHSmqPED3WoiW6hHvsUCTAen1655B9UPAZ3MfjFWUlIxRgWDyd
ubkaalahQ3BgJlKlGBzFjtQTzkP3kI0y+J6N002KfLzVEyNUYucJKZSw/16UHL5PQ6BAuReMCOtU
aUYwvjjT5VxnNsJDoBZdEe4xZO+08z8+xNRliMYpebTlZb9v2tmWeZW2FhDwtUAY6qBPFkV3HNCr
fa6RsEE9rECj3bC+c02QcEX4zxJQW3Bc2tI6j1EhWo+Gg4dPd/LBC3yfMNfNQ/AvzYALCvaMi8I3
jL8LBLOGKMUBMxXslx//Yb2u/zw17zwRtcIAXko5ie1qg+4RZ6+iROfzWBcPAaeZWP3pPjvZF7bv
EDIBZhZXfSNeCI/o+HHWJcnz1qFznIQ0rWHVhOYRUIZS1uAGAkDN9jb17DuD04/8PKvRw6rE1rag
2CJzFuW5UUvVfu3zrGZNmh7MfrO4TcEJtlLViNjCGo/u8WAqXMwjvf7SUZWa2bqTIy2pjSR8AS77
Dv0mmTX3fCEhfeYaSVXPal/ITXpqDPi37QGCjPbtvZNthkLsltRAjuwJbDXsV9NOYGSi331UMEDJ
OZ8A3BnMT/BdwyadDW3xhFyIki9ftD3DxwtZUG22bO6mJ8v7wHcoaJJThXRHjtQLbm/mBJAS0wsI
waSkX6UpLd2brWdbtOGOIWrdEz64YNyTY25sVjzi6yKFfDFHj/2dxB+ssBo087HwQwMyV8dA+YFH
7RDgU0AseJuPAxH23qP+JAtQa33B0uq/yacojfltRkE7ss8NU1Iv6TKQRm25Ov562XU4WHOx03RR
4EX+z+ojHoQJh1Y9/Ya7duVFdO2AfS2mEDMLQoWxZjE7rN9x1QRj885tv7Y+Mg/7Wwc5aAWRlwkF
newOkM9wtUzs1xGxcNBdKsKoTwHS+ws3l/SKE3OCFP6VmxVGgA0BYw9NvGhhQrDfMMYJ8Czl2fsq
u7PLSril+8lB9X9pckdTv3Nh8eYN+WJqtMWHsfrJgHngiVAR7XxeXC/dsAPoPd7pmQsqEglhdog=
`pragma protect end_protected
