   wire                  c0_ddr4_app_correct_en_i;
   wire  [51:0]          c0_ddr4_ecc_err_addr;
   wire  [7:0]           c0_ddr4_ecc_single;
   wire  [7:0]           c0_ddr4_ecc_multiple;

   wire  [27:0]          c0_ddr4_app_addr;
   wire  [2:0]           c0_ddr4_app_cmd;
   wire                  c0_ddr4_app_en;
   wire                  c0_ddr4_app_hi_pri;
   wire  [511:0]         c0_ddr4_app_wdf_data;
   wire                  c0_ddr4_app_wdf_end;
   wire  [63:0]          c0_ddr4_app_wdf_mask;
   wire                  c0_ddr4_app_wdf_wren;
   wire [511:0]          c0_ddr4_app_rd_data;
   wire                  c0_ddr4_app_rd_data_end;
   wire                  c0_ddr4_app_rd_data_valid;
   wire                  c0_ddr4_app_rdy;
   wire                  c0_ddr4_app_wdf_rdy;
   wire                  c0_dbg_clk;
   wire [511:0]          c0_dbg_bus;

   wire                  c1_ddr4_app_correct_en_i;
   wire  [51:0]          c1_ddr4_ecc_err_addr;
   wire  [7:0]           c1_ddr4_ecc_single;
   wire  [7:0]           c1_ddr4_ecc_multiple;

   wire  [27:0]          c1_ddr4_app_addr;
   wire  [2:0]           c1_ddr4_app_cmd;
   wire                  c1_ddr4_app_en;
   wire                  c1_ddr4_app_hi_pri;
   wire  [511:0]         c1_ddr4_app_wdf_data;
   wire                  c1_ddr4_app_wdf_end;
   wire  [63:0]          c1_ddr4_app_wdf_mask;
   wire                  c1_ddr4_app_wdf_wren;
   wire [511:0]          c1_ddr4_app_rd_data;
   wire                  c1_ddr4_app_rd_data_end;
   wire                  c1_ddr4_app_rd_data_valid;
   wire                  c1_ddr4_app_rdy;
   wire                  c1_ddr4_app_wdf_rdy;
   wire                  c1_dbg_clk;
   wire [511:0]          c1_dbg_bus;

   wire                  c2_ddr4_app_correct_en_i;
   wire  [51:0]          c2_ddr4_ecc_err_addr;
   wire  [7:0]           c2_ddr4_ecc_single;
   wire  [7:0]           c2_ddr4_ecc_multiple;

   wire  [27:0]          c2_ddr4_app_addr;
   wire  [2:0]           c2_ddr4_app_cmd;
   wire                  c2_ddr4_app_en;
   wire                  c2_ddr4_app_hi_pri;
   wire  [511:0]         c2_ddr4_app_wdf_data;
   wire                  c2_ddr4_app_wdf_end;
   wire  [63:0]          c2_ddr4_app_wdf_mask;
   wire                  c2_ddr4_app_wdf_wren;
   wire [511:0]          c2_ddr4_app_rd_data;
   wire                  c2_ddr4_app_rd_data_end;
   wire                  c2_ddr4_app_rd_data_valid;
   wire                  c2_ddr4_app_rdy;
   wire                  c2_ddr4_app_wdf_rdy;
   wire                  c2_dbg_clk;
   wire [511:0]          c2_dbg_bus;

   wire                  c3_ddr4_app_correct_en_i;
   wire  [51:0]          c3_ddr4_ecc_err_addr;
   wire  [7:0]           c3_ddr4_ecc_single;
   wire  [7:0]           c3_ddr4_ecc_multiple;

   wire  [27:0]          c3_ddr4_app_addr;
   wire  [2:0]           c3_ddr4_app_cmd;
   wire                  c3_ddr4_app_en;
   wire                  c3_ddr4_app_hi_pri;
   wire  [511:0]         c3_ddr4_app_wdf_data;
   wire                  c3_ddr4_app_wdf_end;
   wire  [63:0]          c3_ddr4_app_wdf_mask;
   wire                  c3_ddr4_app_wdf_wren;
   wire [511:0]          c3_ddr4_app_rd_data;
   wire                  c3_ddr4_app_rd_data_end;
   wire                  c3_ddr4_app_rd_data_valid;
   wire                  c3_ddr4_app_rdy;
   wire                  c3_ddr4_app_wdf_rdy;
   wire                  c3_dbg_clk;
   wire [511:0]          c3_dbg_bus;

